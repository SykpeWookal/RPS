module rpu_thread_control(
  input         clock,
  input         reset,
  input         io_data_stall,
  input         io_control_stall,
  input         io_tkend,
  input         io_addtk,
  input  [31:0] io_time,
  input  [31:0] io_tid,
  input  [31:0] io_ti,
  output        io_wb_pc,
  output        io_pc_we,
  output        io_ifid_clear,
  output        io_ifid_we,
  output        io_idex_clear,
  output        io_idex_we,
  output        io_exmm_clear,
  output        io_exmm_we,
  output        io_mmwb_clear,
  output        io_mmwb_we,
  output        io_thread_id_we,
  output        io_thread_id_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] tt_queue [0:15]; // @[rpu_thread_control.scala 39:21]
  wire  tt_queue_MPORT_1_en; // @[rpu_thread_control.scala 39:21]
  wire [3:0] tt_queue_MPORT_1_addr; // @[rpu_thread_control.scala 39:21]
  wire [63:0] tt_queue_MPORT_1_data; // @[rpu_thread_control.scala 39:21]
  wire  tt_queue_io_thread_id_wdata_MPORT_en; // @[rpu_thread_control.scala 39:21]
  wire [3:0] tt_queue_io_thread_id_wdata_MPORT_addr; // @[rpu_thread_control.scala 39:21]
  wire [63:0] tt_queue_io_thread_id_wdata_MPORT_data; // @[rpu_thread_control.scala 39:21]
  wire [63:0] tt_queue_MPORT_data; // @[rpu_thread_control.scala 39:21]
  wire [3:0] tt_queue_MPORT_addr; // @[rpu_thread_control.scala 39:21]
  wire  tt_queue_MPORT_mask; // @[rpu_thread_control.scala 39:21]
  wire  tt_queue_MPORT_en; // @[rpu_thread_control.scala 39:21]
  reg [3:0] tt_start; // @[rpu_thread_control.scala 40:25]
  reg [3:0] tt_end; // @[rpu_thread_control.scala 41:23]
  reg [1:0] state; // @[rpu_thread_control.scala 44:22]
  wire [3:0] _T_1 = tt_end + 4'h1; // @[rpu_thread_control.scala 49:28]
  wire  _T_2 = _T_1 != tt_start; // @[rpu_thread_control.scala 49:34]
  wire [4:0] _GEN_1 = {{1'd0}, _T_1}; // @[rpu_thread_control.scala 51:30]
  wire [4:0] _GEN_2 = _GEN_1 % 5'h10; // @[rpu_thread_control.scala 51:30]
  wire  _T_5 = state == 2'h3; // @[rpu_thread_control.scala 52:22]
  wire  _T_6 = tt_start != tt_end; // @[rpu_thread_control.scala 52:42]
  wire [3:0] _tt_start_T_1 = tt_start + 4'h1; // @[rpu_thread_control.scala 53:27]
  wire [4:0] _GEN_3 = {{1'd0}, _tt_start_T_1}; // @[rpu_thread_control.scala 53:34]
  wire [4:0] _GEN_4 = _GEN_3 % 5'h10; // @[rpu_thread_control.scala 53:34]
  wire  _T_8 = 2'h0 == state; // @[rpu_thread_control.scala 57:18]
  wire  _GEN_13 = io_tkend ? 1'h0 : 1'h1; // @[rpu_thread_control.scala 39:21 59:23 62:51]
  wire [1:0] _GEN_14 = 2'h3 == state ? 2'h0 : state; // @[rpu_thread_control.scala 57:18 75:13 44:22]
  wire  _T_17 = state == 2'h2; // @[rpu_thread_control.scala 92:22]
  wire  _T_18 = state == 2'h1; // @[rpu_thread_control.scala 105:22]
  wire  _io_pc_we_T = ~io_data_stall; // @[rpu_thread_control.scala 133:17]
  wire  _GEN_23 = io_control_stall | ~io_data_stall; // @[rpu_thread_control.scala 118:34 120:14 133:14]
  wire  _GEN_25 = io_control_stall ? 1'h0 : _io_pc_we_T; // @[rpu_thread_control.scala 118:34 122:16 135:16]
  wire  _GEN_26 = io_control_stall | io_data_stall; // @[rpu_thread_control.scala 118:34 123:19 136:19]
  wire  _GEN_27 = io_control_stall ? 1'h0 : 1'h1; // @[rpu_thread_control.scala 118:34 124:16 137:16]
  wire  _GEN_30 = state == 2'h1 ? 1'h0 : _GEN_23; // @[rpu_thread_control.scala 105:36 107:14]
  wire  _GEN_31 = state == 2'h1 | io_control_stall; // @[rpu_thread_control.scala 105:36 108:19]
  wire  _GEN_32 = state == 2'h1 ? 1'h0 : _GEN_25; // @[rpu_thread_control.scala 105:36 109:16]
  wire  _GEN_33 = state == 2'h1 | _GEN_26; // @[rpu_thread_control.scala 105:36 110:19]
  wire  _GEN_34 = state == 2'h1 ? 1'h0 : _GEN_27; // @[rpu_thread_control.scala 105:36 111:16]
  wire  _GEN_35 = state == 2'h1 ? 1'h0 : 1'h1; // @[rpu_thread_control.scala 105:36 113:16]
  wire  _GEN_38 = state == 2'h2 ? 1'h0 : _T_18; // @[rpu_thread_control.scala 92:35 93:14]
  wire  _GEN_39 = state == 2'h2 ? 1'h0 : _GEN_30; // @[rpu_thread_control.scala 92:35 94:14]
  wire  _GEN_40 = state == 2'h2 ? 1'h0 : _GEN_31; // @[rpu_thread_control.scala 92:35 95:19]
  wire  _GEN_41 = state == 2'h2 ? 1'h0 : _GEN_32; // @[rpu_thread_control.scala 92:35 96:16]
  wire  _GEN_42 = state == 2'h2 ? 1'h0 : _GEN_33; // @[rpu_thread_control.scala 92:35 97:19]
  wire  _GEN_43 = state == 2'h2 ? 1'h0 : _GEN_34; // @[rpu_thread_control.scala 92:35 98:16]
  wire  _GEN_44 = state == 2'h2 ? 1'h0 : _GEN_35; // @[rpu_thread_control.scala 100:16 92:35]
  wire  _GEN_46 = state == 2'h2 ? 1'h0 : 1'h1; // @[rpu_thread_control.scala 102:16 92:35]
  wire [31:0] _GEN_61 = _T_5 ? tt_queue_io_thread_id_wdata_MPORT_data[31:0] : 32'h0; // @[rpu_thread_control.scala 79:24 91:24]
  assign tt_queue_MPORT_1_en = _T_8 & _GEN_13;
  assign tt_queue_MPORT_1_addr = tt_start;
  assign tt_queue_MPORT_1_data = tt_queue[tt_queue_MPORT_1_addr]; // @[rpu_thread_control.scala 39:21]
  assign tt_queue_io_thread_id_wdata_MPORT_en = state == 2'h3;
  assign tt_queue_io_thread_id_wdata_MPORT_addr = tt_start;
  assign tt_queue_io_thread_id_wdata_MPORT_data = tt_queue[tt_queue_io_thread_id_wdata_MPORT_addr]; // @[rpu_thread_control.scala 39:21]
  assign tt_queue_MPORT_data = {io_time,io_tid};
  assign tt_queue_MPORT_addr = tt_end;
  assign tt_queue_MPORT_mask = 1'h1;
  assign tt_queue_MPORT_en = io_addtk & _T_2;
  assign io_wb_pc = _T_5 ? 1'h0 : _GEN_38; // @[rpu_thread_control.scala 79:24 80:14]
  assign io_pc_we = _T_5 ? 1'h0 : _GEN_39; // @[rpu_thread_control.scala 79:24 81:14]
  assign io_ifid_clear = _T_5 ? 1'h0 : _GEN_40; // @[rpu_thread_control.scala 79:24 82:19]
  assign io_ifid_we = _T_5 ? 1'h0 : _GEN_41; // @[rpu_thread_control.scala 79:24 83:16]
  assign io_idex_clear = _T_5 ? 1'h0 : _GEN_42; // @[rpu_thread_control.scala 79:24 84:19]
  assign io_idex_we = _T_5 ? 1'h0 : _GEN_43; // @[rpu_thread_control.scala 79:24 85:16]
  assign io_exmm_clear = _T_5 ? 1'h0 : _GEN_38; // @[rpu_thread_control.scala 79:24 80:14]
  assign io_exmm_we = _T_5 ? 1'h0 : _GEN_44; // @[rpu_thread_control.scala 79:24 87:16]
  assign io_mmwb_clear = _T_5 ? 1'h0 : _T_17; // @[rpu_thread_control.scala 79:24 88:19]
  assign io_mmwb_we = _T_5 ? 1'h0 : _GEN_46; // @[rpu_thread_control.scala 79:24 89:16]
  assign io_thread_id_we = state == 2'h3; // @[rpu_thread_control.scala 79:15]
  assign io_thread_id_wdata = _GEN_61[0];
  always @(posedge clock) begin
    if (tt_queue_MPORT_en & tt_queue_MPORT_mask) begin
      tt_queue[tt_queue_MPORT_addr] <= tt_queue_MPORT_data; // @[rpu_thread_control.scala 39:21]
    end
    if (reset) begin // @[rpu_thread_control.scala 40:25]
      tt_start <= 4'h0; // @[rpu_thread_control.scala 40:25]
    end else if (!(io_addtk & _T_1 != tt_start)) begin // @[rpu_thread_control.scala 49:48]
      if (state == 2'h3 & tt_start != tt_end) begin // @[rpu_thread_control.scala 52:54]
        tt_start <= _GEN_4[3:0]; // @[rpu_thread_control.scala 53:14]
      end
    end
    if (reset) begin // @[rpu_thread_control.scala 41:23]
      tt_end <= 4'h0; // @[rpu_thread_control.scala 41:23]
    end else if (io_addtk & _T_1 != tt_start) begin // @[rpu_thread_control.scala 49:48]
      tt_end <= _GEN_2[3:0]; // @[rpu_thread_control.scala 51:12]
    end
    if (reset) begin // @[rpu_thread_control.scala 44:22]
      state <= 2'h0; // @[rpu_thread_control.scala 44:22]
    end else if (2'h0 == state) begin // @[rpu_thread_control.scala 57:18]
      if (io_tkend) begin // @[rpu_thread_control.scala 59:23]
        state <= 2'h1; // @[rpu_thread_control.scala 61:15]
      end else if (_T_6 & tt_queue_MPORT_1_data[63:32] < io_ti) begin // @[rpu_thread_control.scala 62:79]
        state <= 2'h1; // @[rpu_thread_control.scala 63:15]
      end else begin
        state <= 2'h0; // @[rpu_thread_control.scala 65:15]
      end
    end else if (2'h1 == state) begin // @[rpu_thread_control.scala 57:18]
      state <= 2'h2; // @[rpu_thread_control.scala 69:13]
    end else if (2'h2 == state) begin // @[rpu_thread_control.scala 57:18]
      state <= 2'h3; // @[rpu_thread_control.scala 72:13]
    end else begin
      state <= _GEN_14;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tt_queue[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tt_start = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  tt_end = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rpu_pc_group(
  input         clock,
  input         reset,
  input  [31:0] io_boot_addr_0,
  input  [31:0] io_boot_addr_1,
  input         io_thread_id_we,
  input         io_thread_id_wdata,
  input         io_npc_we,
  input  [31:0] io_npc_wdata,
  output [31:0] io_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc_group_0; // @[rpu_pc_group.scala 25:25]
  reg [31:0] pc_group_1; // @[rpu_pc_group.scala 25:25]
  reg  thread_id; // @[rpu_pc_group.scala 27:22]
  assign io_pc = thread_id ? pc_group_1 : pc_group_0; // @[rpu_pc_group.scala 34:{9,9}]
  always @(posedge clock) begin
    if (reset) begin // @[rpu_pc_group.scala 25:25]
      pc_group_0 <= io_boot_addr_0; // @[rpu_pc_group.scala 25:25]
    end else if (!(io_thread_id_we)) begin // @[rpu_pc_group.scala 29:65]
      if (io_npc_we) begin // @[rpu_pc_group.scala 31:26]
        if (~thread_id) begin // @[rpu_pc_group.scala 32:27]
          pc_group_0 <= io_npc_wdata; // @[rpu_pc_group.scala 32:27]
        end
      end
    end
    if (reset) begin // @[rpu_pc_group.scala 25:25]
      pc_group_1 <= io_boot_addr_1; // @[rpu_pc_group.scala 25:25]
    end else if (!(io_thread_id_we)) begin // @[rpu_pc_group.scala 29:65]
      if (io_npc_we) begin // @[rpu_pc_group.scala 31:26]
        if (thread_id) begin // @[rpu_pc_group.scala 32:27]
          pc_group_1 <= io_npc_wdata; // @[rpu_pc_group.scala 32:27]
        end
      end
    end
    if (io_thread_id_we) begin // @[rpu_pc_group.scala 29:65]
      thread_id <= io_thread_id_wdata; // @[rpu_pc_group.scala 30:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_group_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pc_group_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  thread_id = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegisterFileGroup(
  input         clock,
  input         reset,
  input         io_TID_Change_En,
  input         io_TID_Changed_ID,
  input  [4:0]  io_Raddr1,
  input  [4:0]  io_Raddr2,
  input  [4:0]  io_Raddr3,
  output [31:0] io_Rdata1,
  output [31:0] io_Rdata2,
  output [31:0] io_Rdata3,
  input         io_Write_En,
  input  [4:0]  io_Waddr,
  input  [31:0] io_Wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  reg  TID; // @[RegisterFileGroup.scala 28:16]
  reg [31:0] RegFileGroup_0; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_1; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_2; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_3; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_4; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_5; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_6; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_7; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_8; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_9; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_10; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_11; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_12; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_13; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_14; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_15; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_16; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_17; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_18; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_19; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_20; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_21; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_22; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_23; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_24; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_25; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_26; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_27; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_28; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_29; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_30; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_31; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_32; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_33; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_34; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_35; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_36; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_37; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_38; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_39; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_40; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_41; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_42; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_43; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_44; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_45; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_46; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_47; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_48; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_49; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_50; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_51; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_52; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_53; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_54; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_55; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_56; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_57; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_58; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_59; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_60; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_61; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_62; // @[RegisterFileGroup.scala 30:29]
  reg [31:0] RegFileGroup_63; // @[RegisterFileGroup.scala 30:29]
  wire [5:0] _T_4 = {TID,io_Waddr}; // @[Cat.scala 31:58]
  wire [5:0] _io_Rdata1_T = {TID,io_Raddr1}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_194 = 6'h1 == _io_Rdata1_T ? RegFileGroup_1 : RegFileGroup_0; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_195 = 6'h2 == _io_Rdata1_T ? RegFileGroup_2 : _GEN_194; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_196 = 6'h3 == _io_Rdata1_T ? RegFileGroup_3 : _GEN_195; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_197 = 6'h4 == _io_Rdata1_T ? RegFileGroup_4 : _GEN_196; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_198 = 6'h5 == _io_Rdata1_T ? RegFileGroup_5 : _GEN_197; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_199 = 6'h6 == _io_Rdata1_T ? RegFileGroup_6 : _GEN_198; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_200 = 6'h7 == _io_Rdata1_T ? RegFileGroup_7 : _GEN_199; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_201 = 6'h8 == _io_Rdata1_T ? RegFileGroup_8 : _GEN_200; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_202 = 6'h9 == _io_Rdata1_T ? RegFileGroup_9 : _GEN_201; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_203 = 6'ha == _io_Rdata1_T ? RegFileGroup_10 : _GEN_202; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_204 = 6'hb == _io_Rdata1_T ? RegFileGroup_11 : _GEN_203; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_205 = 6'hc == _io_Rdata1_T ? RegFileGroup_12 : _GEN_204; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_206 = 6'hd == _io_Rdata1_T ? RegFileGroup_13 : _GEN_205; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_207 = 6'he == _io_Rdata1_T ? RegFileGroup_14 : _GEN_206; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_208 = 6'hf == _io_Rdata1_T ? RegFileGroup_15 : _GEN_207; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_209 = 6'h10 == _io_Rdata1_T ? RegFileGroup_16 : _GEN_208; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_210 = 6'h11 == _io_Rdata1_T ? RegFileGroup_17 : _GEN_209; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_211 = 6'h12 == _io_Rdata1_T ? RegFileGroup_18 : _GEN_210; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_212 = 6'h13 == _io_Rdata1_T ? RegFileGroup_19 : _GEN_211; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_213 = 6'h14 == _io_Rdata1_T ? RegFileGroup_20 : _GEN_212; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_214 = 6'h15 == _io_Rdata1_T ? RegFileGroup_21 : _GEN_213; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_215 = 6'h16 == _io_Rdata1_T ? RegFileGroup_22 : _GEN_214; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_216 = 6'h17 == _io_Rdata1_T ? RegFileGroup_23 : _GEN_215; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_217 = 6'h18 == _io_Rdata1_T ? RegFileGroup_24 : _GEN_216; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_218 = 6'h19 == _io_Rdata1_T ? RegFileGroup_25 : _GEN_217; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_219 = 6'h1a == _io_Rdata1_T ? RegFileGroup_26 : _GEN_218; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_220 = 6'h1b == _io_Rdata1_T ? RegFileGroup_27 : _GEN_219; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_221 = 6'h1c == _io_Rdata1_T ? RegFileGroup_28 : _GEN_220; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_222 = 6'h1d == _io_Rdata1_T ? RegFileGroup_29 : _GEN_221; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_223 = 6'h1e == _io_Rdata1_T ? RegFileGroup_30 : _GEN_222; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_224 = 6'h1f == _io_Rdata1_T ? RegFileGroup_31 : _GEN_223; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_225 = 6'h20 == _io_Rdata1_T ? RegFileGroup_32 : _GEN_224; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_226 = 6'h21 == _io_Rdata1_T ? RegFileGroup_33 : _GEN_225; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_227 = 6'h22 == _io_Rdata1_T ? RegFileGroup_34 : _GEN_226; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_228 = 6'h23 == _io_Rdata1_T ? RegFileGroup_35 : _GEN_227; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_229 = 6'h24 == _io_Rdata1_T ? RegFileGroup_36 : _GEN_228; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_230 = 6'h25 == _io_Rdata1_T ? RegFileGroup_37 : _GEN_229; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_231 = 6'h26 == _io_Rdata1_T ? RegFileGroup_38 : _GEN_230; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_232 = 6'h27 == _io_Rdata1_T ? RegFileGroup_39 : _GEN_231; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_233 = 6'h28 == _io_Rdata1_T ? RegFileGroup_40 : _GEN_232; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_234 = 6'h29 == _io_Rdata1_T ? RegFileGroup_41 : _GEN_233; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_235 = 6'h2a == _io_Rdata1_T ? RegFileGroup_42 : _GEN_234; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_236 = 6'h2b == _io_Rdata1_T ? RegFileGroup_43 : _GEN_235; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_237 = 6'h2c == _io_Rdata1_T ? RegFileGroup_44 : _GEN_236; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_238 = 6'h2d == _io_Rdata1_T ? RegFileGroup_45 : _GEN_237; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_239 = 6'h2e == _io_Rdata1_T ? RegFileGroup_46 : _GEN_238; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_240 = 6'h2f == _io_Rdata1_T ? RegFileGroup_47 : _GEN_239; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_241 = 6'h30 == _io_Rdata1_T ? RegFileGroup_48 : _GEN_240; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_242 = 6'h31 == _io_Rdata1_T ? RegFileGroup_49 : _GEN_241; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_243 = 6'h32 == _io_Rdata1_T ? RegFileGroup_50 : _GEN_242; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_244 = 6'h33 == _io_Rdata1_T ? RegFileGroup_51 : _GEN_243; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_245 = 6'h34 == _io_Rdata1_T ? RegFileGroup_52 : _GEN_244; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_246 = 6'h35 == _io_Rdata1_T ? RegFileGroup_53 : _GEN_245; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_247 = 6'h36 == _io_Rdata1_T ? RegFileGroup_54 : _GEN_246; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_248 = 6'h37 == _io_Rdata1_T ? RegFileGroup_55 : _GEN_247; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_249 = 6'h38 == _io_Rdata1_T ? RegFileGroup_56 : _GEN_248; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_250 = 6'h39 == _io_Rdata1_T ? RegFileGroup_57 : _GEN_249; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_251 = 6'h3a == _io_Rdata1_T ? RegFileGroup_58 : _GEN_250; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_252 = 6'h3b == _io_Rdata1_T ? RegFileGroup_59 : _GEN_251; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_253 = 6'h3c == _io_Rdata1_T ? RegFileGroup_60 : _GEN_252; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_254 = 6'h3d == _io_Rdata1_T ? RegFileGroup_61 : _GEN_253; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [31:0] _GEN_255 = 6'h3e == _io_Rdata1_T ? RegFileGroup_62 : _GEN_254; // @[RegisterFileGroup.scala 39:{13,13}]
  wire [5:0] _io_Rdata2_T = {TID,io_Raddr2}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_258 = 6'h1 == _io_Rdata2_T ? RegFileGroup_1 : RegFileGroup_0; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_259 = 6'h2 == _io_Rdata2_T ? RegFileGroup_2 : _GEN_258; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_260 = 6'h3 == _io_Rdata2_T ? RegFileGroup_3 : _GEN_259; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_261 = 6'h4 == _io_Rdata2_T ? RegFileGroup_4 : _GEN_260; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_262 = 6'h5 == _io_Rdata2_T ? RegFileGroup_5 : _GEN_261; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_263 = 6'h6 == _io_Rdata2_T ? RegFileGroup_6 : _GEN_262; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_264 = 6'h7 == _io_Rdata2_T ? RegFileGroup_7 : _GEN_263; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_265 = 6'h8 == _io_Rdata2_T ? RegFileGroup_8 : _GEN_264; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_266 = 6'h9 == _io_Rdata2_T ? RegFileGroup_9 : _GEN_265; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_267 = 6'ha == _io_Rdata2_T ? RegFileGroup_10 : _GEN_266; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_268 = 6'hb == _io_Rdata2_T ? RegFileGroup_11 : _GEN_267; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_269 = 6'hc == _io_Rdata2_T ? RegFileGroup_12 : _GEN_268; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_270 = 6'hd == _io_Rdata2_T ? RegFileGroup_13 : _GEN_269; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_271 = 6'he == _io_Rdata2_T ? RegFileGroup_14 : _GEN_270; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_272 = 6'hf == _io_Rdata2_T ? RegFileGroup_15 : _GEN_271; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_273 = 6'h10 == _io_Rdata2_T ? RegFileGroup_16 : _GEN_272; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_274 = 6'h11 == _io_Rdata2_T ? RegFileGroup_17 : _GEN_273; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_275 = 6'h12 == _io_Rdata2_T ? RegFileGroup_18 : _GEN_274; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_276 = 6'h13 == _io_Rdata2_T ? RegFileGroup_19 : _GEN_275; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_277 = 6'h14 == _io_Rdata2_T ? RegFileGroup_20 : _GEN_276; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_278 = 6'h15 == _io_Rdata2_T ? RegFileGroup_21 : _GEN_277; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_279 = 6'h16 == _io_Rdata2_T ? RegFileGroup_22 : _GEN_278; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_280 = 6'h17 == _io_Rdata2_T ? RegFileGroup_23 : _GEN_279; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_281 = 6'h18 == _io_Rdata2_T ? RegFileGroup_24 : _GEN_280; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_282 = 6'h19 == _io_Rdata2_T ? RegFileGroup_25 : _GEN_281; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_283 = 6'h1a == _io_Rdata2_T ? RegFileGroup_26 : _GEN_282; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_284 = 6'h1b == _io_Rdata2_T ? RegFileGroup_27 : _GEN_283; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_285 = 6'h1c == _io_Rdata2_T ? RegFileGroup_28 : _GEN_284; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_286 = 6'h1d == _io_Rdata2_T ? RegFileGroup_29 : _GEN_285; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_287 = 6'h1e == _io_Rdata2_T ? RegFileGroup_30 : _GEN_286; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_288 = 6'h1f == _io_Rdata2_T ? RegFileGroup_31 : _GEN_287; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_289 = 6'h20 == _io_Rdata2_T ? RegFileGroup_32 : _GEN_288; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_290 = 6'h21 == _io_Rdata2_T ? RegFileGroup_33 : _GEN_289; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_291 = 6'h22 == _io_Rdata2_T ? RegFileGroup_34 : _GEN_290; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_292 = 6'h23 == _io_Rdata2_T ? RegFileGroup_35 : _GEN_291; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_293 = 6'h24 == _io_Rdata2_T ? RegFileGroup_36 : _GEN_292; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_294 = 6'h25 == _io_Rdata2_T ? RegFileGroup_37 : _GEN_293; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_295 = 6'h26 == _io_Rdata2_T ? RegFileGroup_38 : _GEN_294; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_296 = 6'h27 == _io_Rdata2_T ? RegFileGroup_39 : _GEN_295; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_297 = 6'h28 == _io_Rdata2_T ? RegFileGroup_40 : _GEN_296; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_298 = 6'h29 == _io_Rdata2_T ? RegFileGroup_41 : _GEN_297; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_299 = 6'h2a == _io_Rdata2_T ? RegFileGroup_42 : _GEN_298; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_300 = 6'h2b == _io_Rdata2_T ? RegFileGroup_43 : _GEN_299; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_301 = 6'h2c == _io_Rdata2_T ? RegFileGroup_44 : _GEN_300; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_302 = 6'h2d == _io_Rdata2_T ? RegFileGroup_45 : _GEN_301; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_303 = 6'h2e == _io_Rdata2_T ? RegFileGroup_46 : _GEN_302; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_304 = 6'h2f == _io_Rdata2_T ? RegFileGroup_47 : _GEN_303; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_305 = 6'h30 == _io_Rdata2_T ? RegFileGroup_48 : _GEN_304; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_306 = 6'h31 == _io_Rdata2_T ? RegFileGroup_49 : _GEN_305; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_307 = 6'h32 == _io_Rdata2_T ? RegFileGroup_50 : _GEN_306; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_308 = 6'h33 == _io_Rdata2_T ? RegFileGroup_51 : _GEN_307; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_309 = 6'h34 == _io_Rdata2_T ? RegFileGroup_52 : _GEN_308; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_310 = 6'h35 == _io_Rdata2_T ? RegFileGroup_53 : _GEN_309; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_311 = 6'h36 == _io_Rdata2_T ? RegFileGroup_54 : _GEN_310; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_312 = 6'h37 == _io_Rdata2_T ? RegFileGroup_55 : _GEN_311; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_313 = 6'h38 == _io_Rdata2_T ? RegFileGroup_56 : _GEN_312; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_314 = 6'h39 == _io_Rdata2_T ? RegFileGroup_57 : _GEN_313; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_315 = 6'h3a == _io_Rdata2_T ? RegFileGroup_58 : _GEN_314; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_316 = 6'h3b == _io_Rdata2_T ? RegFileGroup_59 : _GEN_315; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_317 = 6'h3c == _io_Rdata2_T ? RegFileGroup_60 : _GEN_316; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_318 = 6'h3d == _io_Rdata2_T ? RegFileGroup_61 : _GEN_317; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [31:0] _GEN_319 = 6'h3e == _io_Rdata2_T ? RegFileGroup_62 : _GEN_318; // @[RegisterFileGroup.scala 40:{13,13}]
  wire [5:0] _io_Rdata3_T = {TID,io_Raddr3}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_322 = 6'h1 == _io_Rdata3_T ? RegFileGroup_1 : RegFileGroup_0; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_323 = 6'h2 == _io_Rdata3_T ? RegFileGroup_2 : _GEN_322; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_324 = 6'h3 == _io_Rdata3_T ? RegFileGroup_3 : _GEN_323; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_325 = 6'h4 == _io_Rdata3_T ? RegFileGroup_4 : _GEN_324; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_326 = 6'h5 == _io_Rdata3_T ? RegFileGroup_5 : _GEN_325; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_327 = 6'h6 == _io_Rdata3_T ? RegFileGroup_6 : _GEN_326; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_328 = 6'h7 == _io_Rdata3_T ? RegFileGroup_7 : _GEN_327; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_329 = 6'h8 == _io_Rdata3_T ? RegFileGroup_8 : _GEN_328; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_330 = 6'h9 == _io_Rdata3_T ? RegFileGroup_9 : _GEN_329; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_331 = 6'ha == _io_Rdata3_T ? RegFileGroup_10 : _GEN_330; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_332 = 6'hb == _io_Rdata3_T ? RegFileGroup_11 : _GEN_331; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_333 = 6'hc == _io_Rdata3_T ? RegFileGroup_12 : _GEN_332; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_334 = 6'hd == _io_Rdata3_T ? RegFileGroup_13 : _GEN_333; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_335 = 6'he == _io_Rdata3_T ? RegFileGroup_14 : _GEN_334; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_336 = 6'hf == _io_Rdata3_T ? RegFileGroup_15 : _GEN_335; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_337 = 6'h10 == _io_Rdata3_T ? RegFileGroup_16 : _GEN_336; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_338 = 6'h11 == _io_Rdata3_T ? RegFileGroup_17 : _GEN_337; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_339 = 6'h12 == _io_Rdata3_T ? RegFileGroup_18 : _GEN_338; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_340 = 6'h13 == _io_Rdata3_T ? RegFileGroup_19 : _GEN_339; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_341 = 6'h14 == _io_Rdata3_T ? RegFileGroup_20 : _GEN_340; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_342 = 6'h15 == _io_Rdata3_T ? RegFileGroup_21 : _GEN_341; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_343 = 6'h16 == _io_Rdata3_T ? RegFileGroup_22 : _GEN_342; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_344 = 6'h17 == _io_Rdata3_T ? RegFileGroup_23 : _GEN_343; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_345 = 6'h18 == _io_Rdata3_T ? RegFileGroup_24 : _GEN_344; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_346 = 6'h19 == _io_Rdata3_T ? RegFileGroup_25 : _GEN_345; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_347 = 6'h1a == _io_Rdata3_T ? RegFileGroup_26 : _GEN_346; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_348 = 6'h1b == _io_Rdata3_T ? RegFileGroup_27 : _GEN_347; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_349 = 6'h1c == _io_Rdata3_T ? RegFileGroup_28 : _GEN_348; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_350 = 6'h1d == _io_Rdata3_T ? RegFileGroup_29 : _GEN_349; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_351 = 6'h1e == _io_Rdata3_T ? RegFileGroup_30 : _GEN_350; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_352 = 6'h1f == _io_Rdata3_T ? RegFileGroup_31 : _GEN_351; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_353 = 6'h20 == _io_Rdata3_T ? RegFileGroup_32 : _GEN_352; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_354 = 6'h21 == _io_Rdata3_T ? RegFileGroup_33 : _GEN_353; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_355 = 6'h22 == _io_Rdata3_T ? RegFileGroup_34 : _GEN_354; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_356 = 6'h23 == _io_Rdata3_T ? RegFileGroup_35 : _GEN_355; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_357 = 6'h24 == _io_Rdata3_T ? RegFileGroup_36 : _GEN_356; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_358 = 6'h25 == _io_Rdata3_T ? RegFileGroup_37 : _GEN_357; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_359 = 6'h26 == _io_Rdata3_T ? RegFileGroup_38 : _GEN_358; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_360 = 6'h27 == _io_Rdata3_T ? RegFileGroup_39 : _GEN_359; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_361 = 6'h28 == _io_Rdata3_T ? RegFileGroup_40 : _GEN_360; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_362 = 6'h29 == _io_Rdata3_T ? RegFileGroup_41 : _GEN_361; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_363 = 6'h2a == _io_Rdata3_T ? RegFileGroup_42 : _GEN_362; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_364 = 6'h2b == _io_Rdata3_T ? RegFileGroup_43 : _GEN_363; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_365 = 6'h2c == _io_Rdata3_T ? RegFileGroup_44 : _GEN_364; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_366 = 6'h2d == _io_Rdata3_T ? RegFileGroup_45 : _GEN_365; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_367 = 6'h2e == _io_Rdata3_T ? RegFileGroup_46 : _GEN_366; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_368 = 6'h2f == _io_Rdata3_T ? RegFileGroup_47 : _GEN_367; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_369 = 6'h30 == _io_Rdata3_T ? RegFileGroup_48 : _GEN_368; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_370 = 6'h31 == _io_Rdata3_T ? RegFileGroup_49 : _GEN_369; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_371 = 6'h32 == _io_Rdata3_T ? RegFileGroup_50 : _GEN_370; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_372 = 6'h33 == _io_Rdata3_T ? RegFileGroup_51 : _GEN_371; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_373 = 6'h34 == _io_Rdata3_T ? RegFileGroup_52 : _GEN_372; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_374 = 6'h35 == _io_Rdata3_T ? RegFileGroup_53 : _GEN_373; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_375 = 6'h36 == _io_Rdata3_T ? RegFileGroup_54 : _GEN_374; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_376 = 6'h37 == _io_Rdata3_T ? RegFileGroup_55 : _GEN_375; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_377 = 6'h38 == _io_Rdata3_T ? RegFileGroup_56 : _GEN_376; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_378 = 6'h39 == _io_Rdata3_T ? RegFileGroup_57 : _GEN_377; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_379 = 6'h3a == _io_Rdata3_T ? RegFileGroup_58 : _GEN_378; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_380 = 6'h3b == _io_Rdata3_T ? RegFileGroup_59 : _GEN_379; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_381 = 6'h3c == _io_Rdata3_T ? RegFileGroup_60 : _GEN_380; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_382 = 6'h3d == _io_Rdata3_T ? RegFileGroup_61 : _GEN_381; // @[RegisterFileGroup.scala 41:{13,13}]
  wire [31:0] _GEN_383 = 6'h3e == _io_Rdata3_T ? RegFileGroup_62 : _GEN_382; // @[RegisterFileGroup.scala 41:{13,13}]
  assign io_Rdata1 = 6'h3f == _io_Rdata1_T ? RegFileGroup_63 : _GEN_255; // @[RegisterFileGroup.scala 39:{13,13}]
  assign io_Rdata2 = 6'h3f == _io_Rdata2_T ? RegFileGroup_63 : _GEN_319; // @[RegisterFileGroup.scala 40:{13,13}]
  assign io_Rdata3 = 6'h3f == _io_Rdata3_T ? RegFileGroup_63 : _GEN_383; // @[RegisterFileGroup.scala 41:{13,13}]
  always @(posedge clock) begin
    if (io_TID_Change_En) begin // @[RegisterFileGroup.scala 33:75]
      TID <= io_TID_Changed_ID; // @[RegisterFileGroup.scala 34:9]
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_0 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h0 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_0 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_1 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_1 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_2 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_2 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_3 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_3 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_4 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h4 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_4 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_5 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h5 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_5 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_6 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h6 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_6 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_7 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h7 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_7 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_8 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h8 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_8 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_9 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h9 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_9 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_10 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'ha == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_10 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_11 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'hb == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_11 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_12 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'hc == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_12 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_13 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'hd == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_13 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_14 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'he == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_14 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_15 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'hf == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_15 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_16 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h10 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_16 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_17 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h11 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_17 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_18 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h12 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_18 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_19 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h13 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_19 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_20 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h14 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_20 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_21 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h15 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_21 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_22 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h16 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_22 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_23 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h17 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_23 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_24 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h18 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_24 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_25 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h19 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_25 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_26 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1a == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_26 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_27 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1b == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_27 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_28 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1c == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_28 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_29 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1d == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_29 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_30 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1e == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_30 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_31 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h1f == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_31 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_32 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h20 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_32 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_33 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h21 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_33 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_34 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h22 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_34 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_35 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h23 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_35 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_36 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h24 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_36 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_37 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h25 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_37 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_38 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h26 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_38 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_39 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h27 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_39 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_40 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h28 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_40 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_41 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h29 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_41 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_42 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2a == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_42 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_43 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2b == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_43 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_44 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2c == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_44 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_45 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2d == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_45 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_46 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2e == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_46 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_47 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h2f == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_47 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_48 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h30 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_48 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_49 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h31 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_49 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_50 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h32 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_50 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_51 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h33 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_51 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_52 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h34 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_52 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_53 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h35 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_53 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_54 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h36 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_54 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_55 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h37 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_55 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_56 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h38 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_56 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_57 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h39 == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_57 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_58 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3a == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_58 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_59 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3b == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_59 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_60 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3c == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_60 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_61 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3d == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_61 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_62 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3e == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_62 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
    if (reset) begin // @[RegisterFileGroup.scala 30:29]
      RegFileGroup_63 <= 32'h0; // @[RegisterFileGroup.scala 30:29]
    end else if (!(io_TID_Change_En)) begin // @[RegisterFileGroup.scala 33:75]
      if (io_Write_En & io_Waddr != 5'h0) begin // @[RegisterFileGroup.scala 35:48]
        if (6'h3f == _T_4) begin // @[RegisterFileGroup.scala 36:38]
          RegFileGroup_63 <= io_Wdata; // @[RegisterFileGroup.scala 36:38]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  TID = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  RegFileGroup_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  RegFileGroup_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  RegFileGroup_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  RegFileGroup_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  RegFileGroup_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  RegFileGroup_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  RegFileGroup_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  RegFileGroup_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  RegFileGroup_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  RegFileGroup_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  RegFileGroup_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  RegFileGroup_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  RegFileGroup_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  RegFileGroup_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  RegFileGroup_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  RegFileGroup_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  RegFileGroup_16 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  RegFileGroup_17 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  RegFileGroup_18 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  RegFileGroup_19 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  RegFileGroup_20 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  RegFileGroup_21 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  RegFileGroup_22 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  RegFileGroup_23 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  RegFileGroup_24 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  RegFileGroup_25 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  RegFileGroup_26 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  RegFileGroup_27 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  RegFileGroup_28 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  RegFileGroup_29 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  RegFileGroup_30 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  RegFileGroup_31 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  RegFileGroup_32 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  RegFileGroup_33 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  RegFileGroup_34 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  RegFileGroup_35 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  RegFileGroup_36 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  RegFileGroup_37 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  RegFileGroup_38 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  RegFileGroup_39 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  RegFileGroup_40 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  RegFileGroup_41 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  RegFileGroup_42 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  RegFileGroup_43 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  RegFileGroup_44 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  RegFileGroup_45 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  RegFileGroup_46 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  RegFileGroup_47 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  RegFileGroup_48 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  RegFileGroup_49 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  RegFileGroup_50 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  RegFileGroup_51 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  RegFileGroup_52 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  RegFileGroup_53 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  RegFileGroup_54 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  RegFileGroup_55 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  RegFileGroup_56 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  RegFileGroup_57 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  RegFileGroup_58 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  RegFileGroup_59 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  RegFileGroup_60 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  RegFileGroup_61 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  RegFileGroup_62 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  RegFileGroup_63 = _RAND_64[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rpu_decoder(
  input  [31:0] io_ir,
  output [5:0]  io_instr_type,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rs3,
  output [4:0]  io_rd,
  output [31:0] io_imm,
  output [11:0] io_CSRAddr
);
  wire  _T_7 = 3'h0 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_8 = 3'h1 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_9 = 3'h2 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_10 = 3'h3 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_11 = 3'h4 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_12 = 3'h5 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_14 = io_ir[31:25] == 7'h0; // @[rpu_decoder.scala 57:31]
  wire  _T_16 = io_ir[31:25] == 7'h20; // @[rpu_decoder.scala 59:38]
  wire [4:0] _GEN_0 = io_ir[31:25] == 7'h20 ? 5'h1b : 5'h0; // @[rpu_decoder.scala 25:17 59:48 60:27]
  wire [4:0] _GEN_1 = io_ir[31:25] == 7'h0 ? 5'h1a : _GEN_0; // @[rpu_decoder.scala 57:40 58:27]
  wire  _T_17 = 3'h6 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire  _T_18 = 3'h7 == io_ir[14:12]; // @[rpu_decoder.scala 40:29]
  wire [4:0] _GEN_2 = 3'h7 == io_ir[14:12] ? 5'h18 : 5'h0; // @[rpu_decoder.scala 25:17 40:29 67:25]
  wire [4:0] _GEN_3 = 3'h6 == io_ir[14:12] ? 5'h17 : _GEN_2; // @[rpu_decoder.scala 40:29 64:25]
  wire [4:0] _GEN_4 = 3'h5 == io_ir[14:12] ? _GEN_1 : _GEN_3; // @[rpu_decoder.scala 40:29]
  wire [4:0] _GEN_5 = 3'h4 == io_ir[14:12] ? 5'h16 : _GEN_4; // @[rpu_decoder.scala 40:29 54:25]
  wire [4:0] _GEN_6 = 3'h3 == io_ir[14:12] ? 5'h15 : _GEN_5; // @[rpu_decoder.scala 40:29 51:25]
  wire [4:0] _GEN_7 = 3'h2 == io_ir[14:12] ? 5'h14 : _GEN_6; // @[rpu_decoder.scala 40:29 48:25]
  wire [4:0] _GEN_8 = 3'h1 == io_ir[14:12] ? 5'h19 : _GEN_7; // @[rpu_decoder.scala 40:29 45:25]
  wire [4:0] _GEN_9 = 3'h0 == io_ir[14:12] ? 5'h13 : _GEN_8; // @[rpu_decoder.scala 40:29 42:25]
  wire [4:0] _GEN_10 = _T_16 ? 5'h1d : 5'h0; // @[rpu_decoder.scala 25:17 76:48 77:27]
  wire [4:0] _GEN_11 = _T_14 ? 5'h1c : _GEN_10; // @[rpu_decoder.scala 74:40 75:27]
  wire [5:0] _GEN_12 = _T_16 ? 6'h23 : 6'h0; // @[rpu_decoder.scala 25:17 95:48 96:27]
  wire [5:0] _GEN_13 = _T_14 ? 6'h22 : _GEN_12; // @[rpu_decoder.scala 93:40 94:27]
  wire [5:0] _GEN_14 = _T_18 ? 6'h25 : 6'h0; // @[rpu_decoder.scala 103:25 25:17 72:29]
  wire [5:0] _GEN_15 = _T_17 ? 6'h24 : _GEN_14; // @[rpu_decoder.scala 100:25 72:29]
  wire [5:0] _GEN_16 = _T_12 ? _GEN_13 : _GEN_15; // @[rpu_decoder.scala 72:29]
  wire [5:0] _GEN_17 = _T_11 ? 6'h21 : _GEN_16; // @[rpu_decoder.scala 72:29 90:25]
  wire [5:0] _GEN_18 = _T_10 ? 6'h20 : _GEN_17; // @[rpu_decoder.scala 72:29 87:25]
  wire [5:0] _GEN_19 = _T_9 ? 6'h1f : _GEN_18; // @[rpu_decoder.scala 72:29 84:25]
  wire [5:0] _GEN_20 = _T_8 ? 6'h1e : _GEN_19; // @[rpu_decoder.scala 72:29 81:25]
  wire [5:0] _GEN_21 = _T_7 ? {{1'd0}, _GEN_11} : _GEN_20; // @[rpu_decoder.scala 72:29]
  wire [3:0] _GEN_22 = _T_12 ? 4'hf : 4'h0; // @[rpu_decoder.scala 108:29 122:25 25:17]
  wire [3:0] _GEN_23 = _T_11 ? 4'he : _GEN_22; // @[rpu_decoder.scala 108:29 119:25]
  wire [3:0] _GEN_24 = _T_9 ? 4'hd : _GEN_23; // @[rpu_decoder.scala 108:29 116:25]
  wire [3:0] _GEN_25 = _T_8 ? 4'hc : _GEN_24; // @[rpu_decoder.scala 108:29 113:25]
  wire [3:0] _GEN_26 = _T_7 ? 4'hb : _GEN_25; // @[rpu_decoder.scala 108:29 110:25]
  wire [4:0] _GEN_27 = _T_9 ? 5'h12 : 5'h0; // @[rpu_decoder.scala 127:29 135:25 25:17]
  wire [4:0] _GEN_28 = _T_8 ? 5'h11 : _GEN_27; // @[rpu_decoder.scala 127:29 132:25]
  wire [4:0] _GEN_29 = _T_7 ? 5'h10 : _GEN_28; // @[rpu_decoder.scala 127:29 129:25]
  wire [3:0] _GEN_30 = _T_18 ? 4'ha : 4'h0; // @[rpu_decoder.scala 140:29 157:25 25:17]
  wire [3:0] _GEN_31 = _T_17 ? 4'h9 : _GEN_30; // @[rpu_decoder.scala 140:29 154:25]
  wire [3:0] _GEN_32 = _T_12 ? 4'h8 : _GEN_31; // @[rpu_decoder.scala 140:29 151:25]
  wire [3:0] _GEN_33 = _T_11 ? 4'h7 : _GEN_32; // @[rpu_decoder.scala 140:29 148:25]
  wire [3:0] _GEN_34 = _T_8 ? 4'h6 : _GEN_33; // @[rpu_decoder.scala 140:29 145:25]
  wire [3:0] _GEN_35 = _T_7 ? 4'h5 : _GEN_34; // @[rpu_decoder.scala 140:29 142:25]
  wire  _T_63 = io_ir[31:25] == 7'h1; // @[rpu_decoder.scala 166:38]
  wire [5:0] _GEN_36 = _T_63 ? 6'h29 : 6'h0; // @[rpu_decoder.scala 170:47 171:27 25:17]
  wire [5:0] _GEN_37 = _T_63 ? 6'h28 : _GEN_36; // @[rpu_decoder.scala 168:47 169:27]
  wire [5:0] _GEN_38 = io_ir[31:25] == 7'h1 ? 6'h27 : _GEN_37; // @[rpu_decoder.scala 166:47 167:27]
  wire [5:0] _GEN_39 = _T_14 ? 6'h26 : _GEN_38; // @[rpu_decoder.scala 164:40 165:27]
  wire [5:0] _GEN_40 = _T_63 ? 6'h2b : 6'h0; // @[rpu_decoder.scala 177:47 178:27 25:17]
  wire [5:0] _GEN_41 = _T_14 ? 6'h2a : _GEN_40; // @[rpu_decoder.scala 175:40 176:27]
  wire [5:0] _GEN_42 = _T_14 ? 6'h2c : 6'h0; // @[rpu_decoder.scala 182:40 183:27 25:17]
  wire [5:0] _GEN_43 = _T_63 ? 6'h2e : 6'h0; // @[rpu_decoder.scala 189:47 190:27 25:17]
  wire [5:0] _GEN_44 = _T_14 ? 6'h2d : _GEN_43; // @[rpu_decoder.scala 187:40 188:27]
  wire [5:0] _GEN_45 = _T_10 ? _GEN_44 : 6'h0; // @[rpu_decoder.scala 162:29 25:17]
  wire [5:0] _GEN_46 = _T_9 ? _GEN_42 : _GEN_45; // @[rpu_decoder.scala 162:29]
  wire [5:0] _GEN_47 = _T_8 ? _GEN_41 : _GEN_46; // @[rpu_decoder.scala 162:29]
  wire [5:0] _GEN_48 = _T_7 ? _GEN_39 : _GEN_47; // @[rpu_decoder.scala 162:29]
  wire [5:0] _GEN_49 = _T_18 ? 6'h34 : 6'h0; // @[rpu_decoder.scala 196:27 219:25 25:17]
  wire [5:0] _GEN_50 = _T_17 ? 6'h33 : _GEN_49; // @[rpu_decoder.scala 196:27 215:25]
  wire [5:0] _GEN_51 = _T_12 ? 6'h32 : _GEN_50; // @[rpu_decoder.scala 196:27 211:25]
  wire [5:0] _GEN_52 = _T_10 ? 6'h31 : _GEN_51; // @[rpu_decoder.scala 196:27 207:25]
  wire [5:0] _GEN_53 = _T_9 ? 6'h30 : _GEN_52; // @[rpu_decoder.scala 196:27 203:25]
  wire [5:0] _GEN_54 = _T_8 ? 6'h2f : _GEN_53; // @[rpu_decoder.scala 196:27 199:25]
  wire [5:0] _GEN_55 = 7'h73 == io_ir[6:0] ? _GEN_54 : 6'h0; // @[rpu_decoder.scala 25:17 26:23]
  wire [5:0] _GEN_56 = 7'hb == io_ir[6:0] ? _GEN_48 : _GEN_55; // @[rpu_decoder.scala 26:23]
  wire [5:0] _GEN_57 = 7'h63 == io_ir[6:0] ? {{2'd0}, _GEN_35} : _GEN_56; // @[rpu_decoder.scala 26:23]
  wire [5:0] _GEN_58 = 7'h23 == io_ir[6:0] ? {{1'd0}, _GEN_29} : _GEN_57; // @[rpu_decoder.scala 26:23]
  wire [5:0] _GEN_59 = 7'h3 == io_ir[6:0] ? {{2'd0}, _GEN_26} : _GEN_58; // @[rpu_decoder.scala 26:23]
  wire [5:0] _GEN_60 = 7'h33 == io_ir[6:0] ? _GEN_21 : _GEN_59; // @[rpu_decoder.scala 26:23]
  wire [5:0] _GEN_61 = 7'h13 == io_ir[6:0] ? {{1'd0}, _GEN_9} : _GEN_60; // @[rpu_decoder.scala 26:23]
  wire [5:0] _GEN_62 = 7'h67 == io_ir[6:0] ? 6'h4 : _GEN_61; // @[rpu_decoder.scala 26:23 37:21]
  wire [5:0] _GEN_63 = 7'h6f == io_ir[6:0] ? 6'h3 : _GEN_62; // @[rpu_decoder.scala 26:23 34:21]
  wire [5:0] _GEN_64 = 7'h17 == io_ir[6:0] ? 6'h2 : _GEN_63; // @[rpu_decoder.scala 26:23 31:21]
  wire  _T_91 = io_instr_type == 6'h2; // @[rpu_decoder.scala 237:23]
  wire  _T_92 = io_instr_type == 6'h1 | _T_91; // @[rpu_decoder.scala 236:42]
  wire [31:0] _io_imm_T = io_ir & 32'hfffff000; // @[rpu_decoder.scala 238:21]
  wire [11:0] _io_imm_T_3 = io_ir[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_imm_T_7 = {_io_imm_T_3,io_ir[19:12],io_ir[20],io_ir[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [20:0] _io_imm_T_10 = io_ir[31] ? 21'h1fffff : 21'h0; // @[Bitwise.scala 74:12]
  wire [32:0] _io_imm_T_12 = {_io_imm_T_10,io_ir[31:20]}; // @[Cat.scala 31:58]
  wire  _T_96 = io_instr_type == 6'h6; // @[rpu_decoder.scala 244:30]
  wire  _T_97 = io_instr_type == 6'h5 | _T_96; // @[rpu_decoder.scala 243:49]
  wire  _T_98 = io_instr_type == 6'h7; // @[rpu_decoder.scala 245:30]
  wire  _T_99 = _T_97 | _T_98; // @[rpu_decoder.scala 244:49]
  wire  _T_100 = io_instr_type == 6'h8; // @[rpu_decoder.scala 246:30]
  wire  _T_101 = _T_99 | _T_100; // @[rpu_decoder.scala 245:49]
  wire  _T_102 = io_instr_type == 6'h9; // @[rpu_decoder.scala 247:30]
  wire  _T_103 = _T_101 | _T_102; // @[rpu_decoder.scala 246:49]
  wire  _T_104 = io_instr_type == 6'ha; // @[rpu_decoder.scala 248:30]
  wire  _T_105 = _T_103 | _T_104; // @[rpu_decoder.scala 247:50]
  wire [19:0] _io_imm_T_15 = io_ir[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_imm_T_19 = {_io_imm_T_15,io_ir[7],io_ir[30:25],io_ir[11:8],1'h0}; // @[Cat.scala 31:58]
  wire  _T_107 = io_instr_type == 6'hc; // @[rpu_decoder.scala 251:30]
  wire  _T_108 = io_instr_type == 6'hb | _T_107; // @[rpu_decoder.scala 250:48]
  wire  _T_109 = io_instr_type == 6'hd; // @[rpu_decoder.scala 252:30]
  wire  _T_110 = _T_108 | _T_109; // @[rpu_decoder.scala 251:48]
  wire  _T_111 = io_instr_type == 6'he; // @[rpu_decoder.scala 253:30]
  wire  _T_112 = _T_110 | _T_111; // @[rpu_decoder.scala 252:48]
  wire  _T_113 = io_instr_type == 6'hf; // @[rpu_decoder.scala 254:30]
  wire  _T_114 = _T_112 | _T_113; // @[rpu_decoder.scala 253:49]
  wire  _T_115 = io_instr_type == 6'h13; // @[rpu_decoder.scala 255:30]
  wire  _T_116 = _T_114 | _T_115; // @[rpu_decoder.scala 254:49]
  wire  _T_117 = io_instr_type == 6'h14; // @[rpu_decoder.scala 256:30]
  wire  _T_118 = _T_116 | _T_117; // @[rpu_decoder.scala 255:50]
  wire  _T_119 = io_instr_type == 6'h15; // @[rpu_decoder.scala 257:30]
  wire  _T_120 = _T_118 | _T_119; // @[rpu_decoder.scala 256:50]
  wire  _T_121 = io_instr_type == 6'h16; // @[rpu_decoder.scala 258:30]
  wire  _T_122 = _T_120 | _T_121; // @[rpu_decoder.scala 257:51]
  wire  _T_123 = io_instr_type == 6'h17; // @[rpu_decoder.scala 259:30]
  wire  _T_124 = _T_122 | _T_123; // @[rpu_decoder.scala 258:50]
  wire  _T_125 = io_instr_type == 6'h18; // @[rpu_decoder.scala 260:30]
  wire  _T_126 = _T_124 | _T_125; // @[rpu_decoder.scala 259:49]
  wire  _T_127 = io_instr_type == 6'h19; // @[rpu_decoder.scala 261:30]
  wire  _T_128 = _T_126 | _T_127; // @[rpu_decoder.scala 260:50]
  wire  _T_129 = io_instr_type == 6'h1a; // @[rpu_decoder.scala 262:30]
  wire  _T_130 = _T_128 | _T_129; // @[rpu_decoder.scala 261:50]
  wire  _T_131 = io_instr_type == 6'h1b; // @[rpu_decoder.scala 263:30]
  wire  _T_132 = _T_130 | _T_131; // @[rpu_decoder.scala 262:50]
  wire [31:0] _io_imm_T_24 = {_io_imm_T_10,io_ir[30:20]}; // @[Cat.scala 31:58]
  wire  _T_134 = io_instr_type == 6'h11; // @[rpu_decoder.scala 266:30]
  wire  _T_135 = io_instr_type == 6'h10 | _T_134; // @[rpu_decoder.scala 265:48]
  wire  _T_136 = io_instr_type == 6'h12; // @[rpu_decoder.scala 267:30]
  wire  _T_137 = _T_135 | _T_136; // @[rpu_decoder.scala 266:48]
  wire [31:0] _io_imm_T_30 = {_io_imm_T_10,io_ir[30:25],io_ir[11:7]}; // @[Cat.scala 31:58]
  wire  _T_139 = io_instr_type == 6'h30; // @[rpu_decoder.scala 270:29]
  wire  _T_140 = io_instr_type == 6'h2f | _T_139; // @[rpu_decoder.scala 269:50]
  wire  _T_141 = io_instr_type == 6'h31; // @[rpu_decoder.scala 271:29]
  wire  _T_142 = _T_140 | _T_141; // @[rpu_decoder.scala 270:50]
  wire  _T_143 = io_instr_type == 6'h32; // @[rpu_decoder.scala 272:29]
  wire  _T_144 = _T_142 | _T_143; // @[rpu_decoder.scala 271:50]
  wire  _T_145 = io_instr_type == 6'h33; // @[rpu_decoder.scala 273:29]
  wire  _T_146 = _T_144 | _T_145; // @[rpu_decoder.scala 272:51]
  wire  _T_147 = io_instr_type == 6'h34; // @[rpu_decoder.scala 274:29]
  wire  _T_148 = _T_146 | _T_147; // @[rpu_decoder.scala 273:51]
  wire [31:0] _io_imm_T_33 = {27'h0,io_ir[19:15]}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_67 = _T_148 ? _io_imm_T_33 : 32'hdeadbeef; // @[rpu_decoder.scala 235:10 274:52 275:12]
  wire [31:0] _GEN_68 = _T_137 ? _io_imm_T_30 : _GEN_67; // @[rpu_decoder.scala 267:49 268:12]
  wire [31:0] _GEN_69 = _T_132 ? _io_imm_T_24 : _GEN_68; // @[rpu_decoder.scala 263:51 264:12]
  wire [31:0] _GEN_70 = _T_105 ? _io_imm_T_19 : _GEN_69; // @[rpu_decoder.scala 248:51 249:12]
  wire [32:0] _GEN_71 = io_instr_type == 6'h4 ? _io_imm_T_12 : {{1'd0}, _GEN_70}; // @[rpu_decoder.scala 241:51 242:12]
  wire [32:0] _GEN_72 = io_instr_type == 6'h3 ? {{1'd0}, _io_imm_T_7} : _GEN_71; // @[rpu_decoder.scala 239:50 240:12]
  wire [32:0] _GEN_73 = _T_92 ? {{1'd0}, _io_imm_T} : _GEN_72; // @[rpu_decoder.scala 237:45 238:12]
  assign io_instr_type = 7'h37 == io_ir[6:0] ? 6'h1 : _GEN_64; // @[rpu_decoder.scala 26:23 28:21]
  assign io_rs1 = io_ir[19:15]; // @[rpu_decoder.scala 226:18]
  assign io_rs2 = io_ir[24:20]; // @[rpu_decoder.scala 227:18]
  assign io_rs3 = io_instr_type == 6'h2b ? io_rd : 5'h0; // @[rpu_decoder.scala 229:45 230:12 232:12]
  assign io_rd = io_ir[11:7]; // @[rpu_decoder.scala 228:17]
  assign io_imm = _GEN_73[31:0];
  assign io_CSRAddr = io_ir[31:20]; // @[rpu_decoder.scala 23:22]
endmodule
module rpu_control(
  input  [5:0] io_instr_type,
  output       io_jump,
  output       io_branch,
  output       io_alu_op1_src,
  output       io_alu_op2_src,
  output [3:0] io_alu_op,
  output [1:0] io_alu_result_src,
  output [2:0] io_comp_op,
  output       io_r2_src,
  output       io_tg_we,
  output       io_ti_we,
  output       io_to,
  output       io_addtk,
  output       io_tkend,
  output       io_mem_write,
  output [3:0] io_mem_op,
  output       io_reg_write,
  output [1:0] io_reg_write_src,
  output [2:0] io_csrType
);
  wire  _T = io_instr_type == 6'h31; // @[rpu_control.scala 31:22]
  wire  _T_1 = io_instr_type == 6'h30; // @[rpu_control.scala 33:28]
  wire  _T_2 = io_instr_type == 6'h2f; // @[rpu_control.scala 35:28]
  wire  _T_3 = io_instr_type == 6'h34; // @[rpu_control.scala 37:28]
  wire  _T_4 = io_instr_type == 6'h33; // @[rpu_control.scala 39:28]
  wire  _T_5 = io_instr_type == 6'h32; // @[rpu_control.scala 41:28]
  wire [2:0] _GEN_0 = io_instr_type == 6'h32 ? 3'h4 : 3'h0; // @[rpu_control.scala 41:50 42:16 44:16]
  wire [2:0] _GEN_1 = io_instr_type == 6'h33 ? 3'h5 : _GEN_0; // @[rpu_control.scala 39:50 40:16]
  wire [2:0] _GEN_2 = io_instr_type == 6'h34 ? 3'h6 : _GEN_1; // @[rpu_control.scala 37:50 38:16]
  wire [2:0] _GEN_3 = io_instr_type == 6'h2f ? 3'h1 : _GEN_2; // @[rpu_control.scala 35:49 36:16]
  wire [2:0] _GEN_4 = io_instr_type == 6'h30 ? 3'h3 : _GEN_3; // @[rpu_control.scala 33:49 34:16]
  wire  _io_jump_T = io_instr_type == 6'h4; // @[rpu_control.scala 47:28]
  wire  _io_jump_T_1 = io_instr_type == 6'h3; // @[rpu_control.scala 47:64]
  wire  _io_jump_T_2 = io_instr_type == 6'h4 | io_instr_type == 6'h3; // @[rpu_control.scala 47:48]
  wire  _io_branch_T = io_instr_type == 6'h5; // @[rpu_control.scala 48:31]
  wire  _io_branch_T_1 = io_instr_type == 6'h6; // @[rpu_control.scala 49:31]
  wire  _io_branch_T_2 = io_instr_type == 6'h5 | _io_branch_T_1; // @[rpu_control.scala 48:50]
  wire  _io_branch_T_3 = io_instr_type == 6'h7; // @[rpu_control.scala 50:31]
  wire  _io_branch_T_4 = _io_branch_T_2 | _io_branch_T_3; // @[rpu_control.scala 49:50]
  wire  _io_branch_T_5 = io_instr_type == 6'h8; // @[rpu_control.scala 51:31]
  wire  _io_branch_T_6 = _io_branch_T_4 | _io_branch_T_5; // @[rpu_control.scala 50:50]
  wire  _io_branch_T_7 = io_instr_type == 6'h9; // @[rpu_control.scala 52:31]
  wire  _io_branch_T_8 = _io_branch_T_6 | _io_branch_T_7; // @[rpu_control.scala 51:50]
  wire  _io_branch_T_9 = io_instr_type == 6'ha; // @[rpu_control.scala 53:31]
  wire  _T_6 = io_instr_type == 6'h2; // @[rpu_control.scala 54:23]
  wire  _T_8 = io_instr_type == 6'h2 | _io_jump_T_1; // @[rpu_control.scala 54:44]
  wire  _T_10 = _T_8 | _io_branch_T; // @[rpu_control.scala 55:42]
  wire  _T_12 = _T_10 | _io_branch_T_1; // @[rpu_control.scala 56:42]
  wire  _T_14 = _T_12 | _io_branch_T_3; // @[rpu_control.scala 57:42]
  wire  _T_16 = _T_14 | _io_branch_T_5; // @[rpu_control.scala 58:42]
  wire  _T_18 = _T_16 | _io_branch_T_7; // @[rpu_control.scala 59:42]
  wire  _T_21 = io_instr_type == 6'h1c; // @[rpu_control.scala 66:23]
  wire  _T_22 = io_instr_type == 6'h1d; // @[rpu_control.scala 67:23]
  wire  _T_23 = io_instr_type == 6'h1c | _T_22; // @[rpu_control.scala 66:42]
  wire  _T_24 = io_instr_type == 6'h1e; // @[rpu_control.scala 68:23]
  wire  _T_25 = _T_23 | _T_24; // @[rpu_control.scala 67:42]
  wire  _T_26 = io_instr_type == 6'h1f; // @[rpu_control.scala 69:23]
  wire  _T_27 = _T_25 | _T_26; // @[rpu_control.scala 68:42]
  wire  _T_28 = io_instr_type == 6'h20; // @[rpu_control.scala 70:23]
  wire  _T_29 = _T_27 | _T_28; // @[rpu_control.scala 69:42]
  wire  _T_30 = io_instr_type == 6'h21; // @[rpu_control.scala 71:23]
  wire  _T_31 = _T_29 | _T_30; // @[rpu_control.scala 70:43]
  wire  _T_32 = io_instr_type == 6'h22; // @[rpu_control.scala 72:23]
  wire  _T_33 = _T_31 | _T_32; // @[rpu_control.scala 71:42]
  wire  _T_34 = io_instr_type == 6'h23; // @[rpu_control.scala 73:23]
  wire  _T_35 = _T_33 | _T_34; // @[rpu_control.scala 72:42]
  wire  _T_36 = io_instr_type == 6'h24; // @[rpu_control.scala 74:23]
  wire  _T_37 = _T_35 | _T_36; // @[rpu_control.scala 73:42]
  wire  _T_39 = _T_37 | _T_21; // @[rpu_control.scala 74:41]
  wire  _T_42 = 6'hb == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_45 = 6'hc == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_48 = 6'hd == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_51 = 6'he == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_54 = 6'hf == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_57 = 6'h10 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_60 = 6'h11 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_63 = 6'h12 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_84 = 6'h5 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_87 = 6'h6 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_90 = 6'h7 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_93 = 6'h8 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_96 = 6'h9 == io_instr_type; // @[rpu_control.scala 82:26]
  wire  _T_99 = 6'ha == io_instr_type; // @[rpu_control.scala 82:26]
  wire [3:0] _GEN_8 = 6'h34 == io_instr_type ? 4'hd : 4'h0; // @[rpu_control.scala 210:17 81:13 82:26]
  wire [3:0] _GEN_9 = 6'h33 == io_instr_type ? 4'hd : _GEN_8; // @[rpu_control.scala 207:17 82:26]
  wire [3:0] _GEN_10 = 6'h32 == io_instr_type ? 4'hd : _GEN_9; // @[rpu_control.scala 204:17 82:26]
  wire [3:0] _GEN_11 = 6'h31 == io_instr_type ? 4'hd : _GEN_10; // @[rpu_control.scala 201:17 82:26]
  wire [3:0] _GEN_12 = 6'h30 == io_instr_type ? 4'hd : _GEN_11; // @[rpu_control.scala 198:17 82:26]
  wire [3:0] _GEN_13 = 6'h2f == io_instr_type ? 4'hd : _GEN_12; // @[rpu_control.scala 195:17 82:26]
  wire [3:0] _GEN_14 = 6'h1b == io_instr_type ? 4'h7 : _GEN_13; // @[rpu_control.scala 192:17 82:26]
  wire [3:0] _GEN_15 = 6'h23 == io_instr_type ? 4'h7 : _GEN_14; // @[rpu_control.scala 189:17 82:26]
  wire [3:0] _GEN_16 = 6'h1a == io_instr_type ? 4'h8 : _GEN_15; // @[rpu_control.scala 186:17 82:26]
  wire [3:0] _GEN_17 = 6'h22 == io_instr_type ? 4'h8 : _GEN_16; // @[rpu_control.scala 183:17 82:26]
  wire [3:0] _GEN_18 = 6'h19 == io_instr_type ? 4'h6 : _GEN_17; // @[rpu_control.scala 180:17 82:26]
  wire [3:0] _GEN_19 = 6'h1e == io_instr_type ? 4'h6 : _GEN_18; // @[rpu_control.scala 177:17 82:26]
  wire [3:0] _GEN_20 = 6'h18 == io_instr_type ? 4'h5 : _GEN_19; // @[rpu_control.scala 174:17 82:26]
  wire [3:0] _GEN_21 = 6'h25 == io_instr_type ? 4'h5 : _GEN_20; // @[rpu_control.scala 171:17 82:26]
  wire [3:0] _GEN_22 = 6'h17 == io_instr_type ? 4'h4 : _GEN_21; // @[rpu_control.scala 168:17 82:26]
  wire [3:0] _GEN_23 = 6'h24 == io_instr_type ? 4'h4 : _GEN_22; // @[rpu_control.scala 165:17 82:26]
  wire [3:0] _GEN_24 = 6'h16 == io_instr_type ? 4'h3 : _GEN_23; // @[rpu_control.scala 162:17 82:26]
  wire [3:0] _GEN_25 = 6'h21 == io_instr_type ? 4'h3 : _GEN_24; // @[rpu_control.scala 159:17 82:26]
  wire [3:0] _GEN_26 = 6'h15 == io_instr_type ? 4'hb : _GEN_25; // @[rpu_control.scala 156:17 82:26]
  wire [3:0] _GEN_27 = 6'h20 == io_instr_type ? 4'hb : _GEN_26; // @[rpu_control.scala 153:17 82:26]
  wire [3:0] _GEN_28 = 6'h14 == io_instr_type ? 4'ha : _GEN_27; // @[rpu_control.scala 150:17 82:26]
  wire [3:0] _GEN_29 = 6'h1f == io_instr_type ? 4'ha : _GEN_28; // @[rpu_control.scala 147:17 82:26]
  wire [3:0] _GEN_30 = 6'h1d == io_instr_type ? 4'h2 : _GEN_29; // @[rpu_control.scala 144:17 82:26]
  wire [3:0] _GEN_31 = 6'ha == io_instr_type ? 4'h1 : _GEN_30; // @[rpu_control.scala 141:17 82:26]
  wire [3:0] _GEN_32 = 6'h9 == io_instr_type ? 4'h1 : _GEN_31; // @[rpu_control.scala 138:17 82:26]
  wire [3:0] _GEN_33 = 6'h8 == io_instr_type ? 4'h1 : _GEN_32; // @[rpu_control.scala 135:17 82:26]
  wire [3:0] _GEN_34 = 6'h7 == io_instr_type ? 4'h1 : _GEN_33; // @[rpu_control.scala 132:17 82:26]
  wire [3:0] _GEN_35 = 6'h6 == io_instr_type ? 4'h1 : _GEN_34; // @[rpu_control.scala 129:17 82:26]
  wire [3:0] _GEN_36 = 6'h5 == io_instr_type ? 4'h1 : _GEN_35; // @[rpu_control.scala 126:17 82:26]
  wire [3:0] _GEN_37 = 6'h13 == io_instr_type ? 4'h1 : _GEN_36; // @[rpu_control.scala 123:17 82:26]
  wire [3:0] _GEN_38 = 6'h1c == io_instr_type ? 4'h1 : _GEN_37; // @[rpu_control.scala 120:17 82:26]
  wire [3:0] _GEN_39 = 6'h2 == io_instr_type ? 4'h1 : _GEN_38; // @[rpu_control.scala 117:17 82:26]
  wire [3:0] _GEN_40 = 6'h4 == io_instr_type ? 4'h1 : _GEN_39; // @[rpu_control.scala 114:17 82:26]
  wire [3:0] _GEN_41 = 6'h3 == io_instr_type ? 4'h1 : _GEN_40; // @[rpu_control.scala 111:17 82:26]
  wire [3:0] _GEN_42 = 6'h1 == io_instr_type ? 4'h9 : _GEN_41; // @[rpu_control.scala 108:17 82:26]
  wire [3:0] _GEN_43 = 6'h12 == io_instr_type ? 4'h1 : _GEN_42; // @[rpu_control.scala 105:17 82:26]
  wire [3:0] _GEN_44 = 6'h11 == io_instr_type ? 4'h1 : _GEN_43; // @[rpu_control.scala 102:17 82:26]
  wire [3:0] _GEN_45 = 6'h10 == io_instr_type ? 4'h1 : _GEN_44; // @[rpu_control.scala 82:26 99:17]
  wire [3:0] _GEN_46 = 6'hf == io_instr_type ? 4'h1 : _GEN_45; // @[rpu_control.scala 82:26 96:17]
  wire [3:0] _GEN_47 = 6'he == io_instr_type ? 4'h1 : _GEN_46; // @[rpu_control.scala 82:26 93:17]
  wire [3:0] _GEN_48 = 6'hd == io_instr_type ? 4'h1 : _GEN_47; // @[rpu_control.scala 82:26 90:17]
  wire [3:0] _GEN_49 = 6'hc == io_instr_type ? 4'h1 : _GEN_48; // @[rpu_control.scala 82:26 87:17]
  wire  _T_169 = io_instr_type == 6'h29; // @[rpu_control.scala 215:23]
  wire  _T_170 = io_instr_type == 6'h28; // @[rpu_control.scala 217:30]
  wire [1:0] _GEN_51 = io_instr_type == 6'h28 ? 2'h2 : 2'h0; // @[rpu_control.scala 217:52 218:23 220:23]
  wire [2:0] _GEN_53 = _T_99 ? 3'h6 : 3'h0; // @[rpu_control.scala 223:14 224:26 241:18]
  wire [2:0] _GEN_54 = _T_96 ? 3'h4 : _GEN_53; // @[rpu_control.scala 224:26 238:18]
  wire [2:0] _GEN_55 = _T_93 ? 3'h5 : _GEN_54; // @[rpu_control.scala 224:26 235:18]
  wire [2:0] _GEN_56 = _T_90 ? 3'h3 : _GEN_55; // @[rpu_control.scala 224:26 232:18]
  wire [2:0] _GEN_57 = _T_87 ? 3'h2 : _GEN_56; // @[rpu_control.scala 224:26 229:18]
  wire  _T_189 = io_instr_type == 6'h2b; // @[rpu_control.scala 245:23]
  wire  _io_to_T = io_instr_type == 6'h2a; // @[rpu_control.scala 252:26]
  wire  _io_to_T_2 = io_instr_type == 6'h2a | _T_189; // @[rpu_control.scala 252:47]
  wire  _io_to_T_3 = io_instr_type == 6'h2c; // @[rpu_control.scala 254:26]
  wire  _io_mem_write_T_1 = io_instr_type == 6'h11; // @[rpu_control.scala 258:33]
  wire  _io_mem_write_T_2 = io_instr_type == 6'h10 | _io_mem_write_T_1; // @[rpu_control.scala 257:51]
  wire  _io_mem_write_T_3 = io_instr_type == 6'h12; // @[rpu_control.scala 259:33]
  wire  _io_mem_write_T_4 = _io_mem_write_T_2 | _io_mem_write_T_3; // @[rpu_control.scala 258:51]
  wire [1:0] _GEN_60 = 6'h2a == io_instr_type ? 2'h3 : 2'h0; // @[rpu_control.scala 261:13 262:26 291:17]
  wire [1:0] _GEN_61 = _T_48 ? 2'h3 : _GEN_60; // @[rpu_control.scala 262:26 288:17]
  wire [2:0] _GEN_62 = _T_54 ? 3'h5 : {{1'd0}, _GEN_61}; // @[rpu_control.scala 262:26 285:17]
  wire [2:0] _GEN_63 = _T_45 ? 3'h2 : _GEN_62; // @[rpu_control.scala 262:26 282:17]
  wire [2:0] _GEN_64 = _T_51 ? 3'h4 : _GEN_63; // @[rpu_control.scala 262:26 279:17]
  wire [2:0] _GEN_65 = _T_42 ? 3'h1 : _GEN_64; // @[rpu_control.scala 262:26 276:17]
  wire [3:0] _GEN_66 = 6'h2b == io_instr_type ? 4'h8 : {{1'd0}, _GEN_65}; // @[rpu_control.scala 262:26 273:17]
  wire [3:0] _GEN_67 = _T_63 ? 4'h8 : _GEN_66; // @[rpu_control.scala 262:26 270:17]
  wire [3:0] _GEN_68 = _T_60 ? 4'h7 : _GEN_67; // @[rpu_control.scala 262:26 267:17]
  wire  _io_reg_write_T_2 = io_instr_type == 6'h1 | _T_6; // @[rpu_control.scala 294:52]
  wire  _io_reg_write_T_3 = io_instr_type == 6'h13; // @[rpu_control.scala 296:33]
  wire  _io_reg_write_T_4 = _io_reg_write_T_2 | _io_reg_write_T_3; // @[rpu_control.scala 295:54]
  wire  _io_reg_write_T_5 = io_instr_type == 6'h14; // @[rpu_control.scala 297:33]
  wire  _io_reg_write_T_6 = _io_reg_write_T_4 | _io_reg_write_T_5; // @[rpu_control.scala 296:53]
  wire  _io_reg_write_T_8 = _io_reg_write_T_6 | _T_28; // @[rpu_control.scala 297:53]
  wire  _io_reg_write_T_9 = io_instr_type == 6'h16; // @[rpu_control.scala 299:33]
  wire  _io_reg_write_T_10 = _io_reg_write_T_8 | _io_reg_write_T_9; // @[rpu_control.scala 298:53]
  wire  _io_reg_write_T_11 = io_instr_type == 6'h17; // @[rpu_control.scala 300:33]
  wire  _io_reg_write_T_12 = _io_reg_write_T_10 | _io_reg_write_T_11; // @[rpu_control.scala 299:53]
  wire  _io_reg_write_T_13 = io_instr_type == 6'h18; // @[rpu_control.scala 301:33]
  wire  _io_reg_write_T_14 = _io_reg_write_T_12 | _io_reg_write_T_13; // @[rpu_control.scala 300:52]
  wire  _io_reg_write_T_15 = io_instr_type == 6'h19; // @[rpu_control.scala 302:33]
  wire  _io_reg_write_T_16 = _io_reg_write_T_14 | _io_reg_write_T_15; // @[rpu_control.scala 301:53]
  wire  _io_reg_write_T_17 = io_instr_type == 6'h1a; // @[rpu_control.scala 303:33]
  wire  _io_reg_write_T_18 = _io_reg_write_T_16 | _io_reg_write_T_17; // @[rpu_control.scala 302:53]
  wire  _io_reg_write_T_19 = io_instr_type == 6'h1b; // @[rpu_control.scala 304:33]
  wire  _io_reg_write_T_20 = _io_reg_write_T_18 | _io_reg_write_T_19; // @[rpu_control.scala 303:53]
  wire  _io_reg_write_T_22 = _io_reg_write_T_20 | _T_21; // @[rpu_control.scala 304:53]
  wire  _io_reg_write_T_24 = _io_reg_write_T_22 | _T_22; // @[rpu_control.scala 305:52]
  wire  _io_reg_write_T_26 = _io_reg_write_T_24 | _T_24; // @[rpu_control.scala 306:52]
  wire  _io_reg_write_T_28 = _io_reg_write_T_26 | _T_26; // @[rpu_control.scala 307:52]
  wire  _io_reg_write_T_30 = _io_reg_write_T_28 | _T_28; // @[rpu_control.scala 308:52]
  wire  _io_reg_write_T_32 = _io_reg_write_T_30 | _T_30; // @[rpu_control.scala 309:53]
  wire  _io_reg_write_T_34 = _io_reg_write_T_32 | _T_32; // @[rpu_control.scala 310:52]
  wire  _io_reg_write_T_36 = _io_reg_write_T_34 | _T_34; // @[rpu_control.scala 311:52]
  wire  _io_reg_write_T_38 = _io_reg_write_T_36 | _T_36; // @[rpu_control.scala 312:52]
  wire  _io_reg_write_T_39 = io_instr_type == 6'h25; // @[rpu_control.scala 314:33]
  wire  _io_reg_write_T_40 = _io_reg_write_T_38 | _io_reg_write_T_39; // @[rpu_control.scala 313:51]
  wire  _io_reg_write_T_41 = io_instr_type == 6'hb; // @[rpu_control.scala 315:33]
  wire  _io_reg_write_T_42 = _io_reg_write_T_40 | _io_reg_write_T_41; // @[rpu_control.scala 314:52]
  wire  _io_reg_write_T_43 = io_instr_type == 6'hc; // @[rpu_control.scala 316:33]
  wire  _io_reg_write_T_44 = _io_reg_write_T_42 | _io_reg_write_T_43; // @[rpu_control.scala 315:51]
  wire  _io_reg_write_T_45 = io_instr_type == 6'hd; // @[rpu_control.scala 317:33]
  wire  _io_reg_write_T_46 = _io_reg_write_T_44 | _io_reg_write_T_45; // @[rpu_control.scala 316:51]
  wire  _io_reg_write_T_47 = io_instr_type == 6'he; // @[rpu_control.scala 318:33]
  wire  _io_reg_write_T_48 = _io_reg_write_T_46 | _io_reg_write_T_47; // @[rpu_control.scala 317:51]
  wire  _io_reg_write_T_49 = io_instr_type == 6'hf; // @[rpu_control.scala 319:33]
  wire  _io_reg_write_T_50 = _io_reg_write_T_48 | _io_reg_write_T_49; // @[rpu_control.scala 318:52]
  wire  _io_reg_write_T_52 = _io_reg_write_T_50 | _io_jump_T; // @[rpu_control.scala 319:52]
  wire  _io_reg_write_T_54 = _io_reg_write_T_52 | _io_jump_T_1; // @[rpu_control.scala 320:53]
  wire  _io_reg_write_T_56 = _io_reg_write_T_54 | _T_170; // @[rpu_control.scala 321:52]
  wire  _io_reg_write_T_58 = _io_reg_write_T_56 | _T_169; // @[rpu_control.scala 322:54]
  wire  _io_reg_write_T_60 = _io_reg_write_T_58 | _io_to_T; // @[rpu_control.scala 323:54]
  wire  _io_reg_write_T_62 = _io_reg_write_T_60 | _T_2; // @[rpu_control.scala 324:54]
  wire  _io_reg_write_T_64 = _io_reg_write_T_62 | _T_1; // @[rpu_control.scala 325:54]
  wire  _io_reg_write_T_66 = _io_reg_write_T_64 | _T; // @[rpu_control.scala 326:54]
  wire  _io_reg_write_T_68 = _io_reg_write_T_66 | _T_5; // @[rpu_control.scala 327:54]
  wire  _io_reg_write_T_70 = _io_reg_write_T_68 | _T_4; // @[rpu_control.scala 328:55]
  wire  _T_222 = _io_reg_write_T_41 | _io_reg_write_T_43; // @[rpu_control.scala 331:41]
  wire  _T_224 = _T_222 | _io_reg_write_T_45; // @[rpu_control.scala 332:41]
  wire  _T_226 = _T_224 | _io_reg_write_T_47; // @[rpu_control.scala 333:41]
  wire  _T_228 = _T_226 | _io_reg_write_T_49; // @[rpu_control.scala 334:42]
  wire  _T_230 = _T_228 | _io_to_T; // @[rpu_control.scala 335:42]
  wire [1:0] _GEN_70 = _io_jump_T_2 ? 2'h2 : 2'h1; // @[rpu_control.scala 339:51 340:22 342:22]
  assign io_jump = io_instr_type == 6'h4 | io_instr_type == 6'h3; // @[rpu_control.scala 47:48]
  assign io_branch = _io_branch_T_8 | _io_branch_T_9; // @[rpu_control.scala 52:51]
  assign io_alu_op1_src = _T_18 | _io_branch_T_9; // @[rpu_control.scala 60:43]
  assign io_alu_op2_src = _T_39 ? 1'h0 : 1'h1; // @[rpu_control.scala 75:43 76:20 78:20]
  assign io_alu_op = 6'hb == io_instr_type ? 4'h1 : _GEN_49; // @[rpu_control.scala 82:26 84:17]
  assign io_alu_result_src = io_instr_type == 6'h29 ? 2'h1 : _GEN_51; // @[rpu_control.scala 215:45 216:23]
  assign io_comp_op = _T_84 ? 3'h1 : _GEN_57; // @[rpu_control.scala 224:26 226:18]
  assign io_r2_src = io_instr_type == 6'h2b; // @[rpu_control.scala 245:23]
  assign io_tg_we = io_instr_type == 6'h26; // @[rpu_control.scala 250:29]
  assign io_ti_we = io_instr_type == 6'h27; // @[rpu_control.scala 251:29]
  assign io_to = _io_to_T_2 | _io_to_T_3; // @[rpu_control.scala 253:47]
  assign io_addtk = io_instr_type == 6'h2e; // @[rpu_control.scala 255:29]
  assign io_tkend = io_instr_type == 6'h2d; // @[rpu_control.scala 256:29]
  assign io_mem_write = _io_mem_write_T_4 | _T_189; // @[rpu_control.scala 259:51]
  assign io_mem_op = _T_57 ? 4'h6 : _GEN_68; // @[rpu_control.scala 262:26 264:17]
  assign io_reg_write = _io_reg_write_T_70 | _T_3; // @[rpu_control.scala 329:55]
  assign io_reg_write_src = _T_230 ? 2'h0 : _GEN_70; // @[rpu_control.scala 336:45 337:22]
  assign io_csrType = io_instr_type == 6'h31 ? 3'h3 : _GEN_4; // @[rpu_control.scala 31:43 32:16]
endmodule
module rpu_alu(
  input  [31:0] io_op_a,
  input  [31:0] io_op_b,
  input  [31:0] io_csrResult,
  input  [3:0]  io_operation,
  output [31:0] io_result
);
  wire [31:0] _io_result_T_1 = io_op_a + io_op_b; // @[rpu_alu.scala 18:28]
  wire [31:0] _io_result_T_3 = io_op_a - io_op_b; // @[rpu_alu.scala 21:28]
  wire [31:0] _io_result_T_4 = io_op_a & io_op_b; // @[rpu_alu.scala 24:28]
  wire [31:0] _io_result_T_5 = io_op_a | io_op_b; // @[rpu_alu.scala 27:28]
  wire [31:0] _io_result_T_6 = io_op_a ^ io_op_b; // @[rpu_alu.scala 30:28]
  wire [62:0] _GEN_13 = {{31'd0}, io_op_a}; // @[rpu_alu.scala 33:28]
  wire [62:0] _io_result_T_8 = _GEN_13 << io_op_b[4:0]; // @[rpu_alu.scala 33:28]
  wire [31:0] _io_result_T_9 = io_op_a; // @[rpu_alu.scala 36:29]
  wire [31:0] _io_result_T_12 = $signed(io_op_a) >>> io_op_b[4:0]; // @[rpu_alu.scala 36:54]
  wire [31:0] _io_result_T_14 = io_op_a >> io_op_b[4:0]; // @[rpu_alu.scala 39:28]
  wire [31:0] _io_result_T_16 = io_op_b; // @[rpu_alu.scala 45:45]
  wire [31:0] _GEN_0 = 4'h0 == io_operation ? 32'hdeadbeef : 32'h0; // @[rpu_alu.scala 15:13 16:24 54:17]
  wire [31:0] _GEN_1 = 4'hd == io_operation ? io_csrResult : _GEN_0; // @[rpu_alu.scala 16:24 51:17]
  wire [31:0] _GEN_2 = 4'hb == io_operation ? {{31'd0}, io_op_a < io_op_b} : _GEN_1; // @[rpu_alu.scala 16:24 48:17]
  wire [31:0] _GEN_3 = 4'ha == io_operation ? {{31'd0}, $signed(_io_result_T_9) < $signed(_io_result_T_16)} : _GEN_2; // @[rpu_alu.scala 16:24 45:17]
  wire [31:0] _GEN_4 = 4'h9 == io_operation ? io_op_b : _GEN_3; // @[rpu_alu.scala 16:24 42:17]
  wire [31:0] _GEN_5 = 4'h8 == io_operation ? _io_result_T_14 : _GEN_4; // @[rpu_alu.scala 16:24 39:17]
  wire [31:0] _GEN_6 = 4'h7 == io_operation ? _io_result_T_12 : _GEN_5; // @[rpu_alu.scala 16:24 36:17]
  wire [62:0] _GEN_7 = 4'h6 == io_operation ? _io_result_T_8 : {{31'd0}, _GEN_6}; // @[rpu_alu.scala 16:24 33:17]
  wire [62:0] _GEN_8 = 4'h3 == io_operation ? {{31'd0}, _io_result_T_6} : _GEN_7; // @[rpu_alu.scala 16:24 30:17]
  wire [62:0] _GEN_9 = 4'h4 == io_operation ? {{31'd0}, _io_result_T_5} : _GEN_8; // @[rpu_alu.scala 16:24 27:17]
  wire [62:0] _GEN_10 = 4'h5 == io_operation ? {{31'd0}, _io_result_T_4} : _GEN_9; // @[rpu_alu.scala 16:24 24:17]
  wire [62:0] _GEN_11 = 4'h2 == io_operation ? {{31'd0}, _io_result_T_3} : _GEN_10; // @[rpu_alu.scala 16:24 21:17]
  wire [62:0] _GEN_12 = 4'h1 == io_operation ? {{31'd0}, _io_result_T_1} : _GEN_11; // @[rpu_alu.scala 16:24 18:17]
  assign io_result = _GEN_12[31:0];
endmodule
module rpu_comp(
  input  [2:0]  io_comp_op,
  input  [31:0] io_op_a,
  input  [31:0] io_op_b,
  output        io_result
);
  wire  _GEN_0 = 3'h6 == io_comp_op & io_op_a >= io_op_b; // @[rpu_alu.scala 67:13 68:22 85:17]
  wire  _GEN_1 = 3'h5 == io_comp_op ? $signed(io_op_a) >= $signed(io_op_b) : _GEN_0; // @[rpu_alu.scala 68:22 82:17]
  wire  _GEN_2 = 3'h4 == io_comp_op ? io_op_a < io_op_b : _GEN_1; // @[rpu_alu.scala 68:22 79:17]
  wire  _GEN_3 = 3'h3 == io_comp_op ? $signed(io_op_a) < $signed(io_op_b) : _GEN_2; // @[rpu_alu.scala 68:22 76:17]
  wire  _GEN_4 = 3'h2 == io_comp_op ? io_op_a != io_op_b : _GEN_3; // @[rpu_alu.scala 68:22 73:17]
  assign io_result = 3'h1 == io_comp_op ? io_op_a == io_op_b : _GEN_4; // @[rpu_alu.scala 68:22 70:17]
endmodule
module rpu_time_unit(
  input         clock,
  input         reset,
  input         io_std_clk,
  input         io_ti_we,
  input  [31:0] io_ti_wdata,
  input         io_tg_we,
  input  [31:0] io_tg_wdata,
  output [31:0] io_ti
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  tick; // @[rpu_time_unit.scala 20:21]
  wire  _GEN_0 = ~io_std_clk ? 1'h0 : tick; // @[rpu_time_unit.scala 23:40 24:10 26:10]
  wire  _GEN_1 = io_std_clk & ~tick | _GEN_0; // @[rpu_time_unit.scala 21:52 22:10]
  reg [31:0] ti; // @[rpu_time_unit.scala 29:19]
  reg [31:0] tg; // @[rpu_time_unit.scala 30:19]
  reg [31:0] cnt; // @[rpu_time_unit.scala 31:20]
  wire [31:0] _cnt_T_1 = cnt + 32'h1; // @[rpu_time_unit.scala 34:16]
  wire [31:0] _ti_T_1 = ti + 32'h1; // @[rpu_time_unit.scala 43:14]
  assign io_ti = ti; // @[rpu_time_unit.scala 54:9]
  always @(posedge clock) begin
    if (reset) begin // @[rpu_time_unit.scala 20:21]
      tick <= 1'h0; // @[rpu_time_unit.scala 20:21]
    end else if (tick) begin // @[rpu_time_unit.scala 33:15]
      tick <= 1'h0; // @[rpu_time_unit.scala 35:10]
    end else begin
      tick <= _GEN_1;
    end
    if (reset) begin // @[rpu_time_unit.scala 29:19]
      ti <= 32'h0; // @[rpu_time_unit.scala 29:19]
    end else if (io_ti_we) begin // @[rpu_time_unit.scala 40:19]
      ti <= io_ti_wdata; // @[rpu_time_unit.scala 41:8]
    end else if (cnt == tg) begin // @[rpu_time_unit.scala 42:28]
      ti <= _ti_T_1; // @[rpu_time_unit.scala 43:8]
    end
    if (reset) begin // @[rpu_time_unit.scala 30:19]
      tg <= 32'h0; // @[rpu_time_unit.scala 30:19]
    end else if (io_tg_we) begin // @[rpu_time_unit.scala 48:19]
      tg <= io_tg_wdata; // @[rpu_time_unit.scala 49:8]
    end
    if (reset) begin // @[rpu_time_unit.scala 31:20]
      cnt <= 32'h0; // @[rpu_time_unit.scala 31:20]
    end else if (tick) begin // @[rpu_time_unit.scala 33:15]
      cnt <= _cnt_T_1; // @[rpu_time_unit.scala 34:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tick = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ti = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  tg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cnt = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [2:0]  io_CSRType,
  input  [11:0] io_CSRAddr,
  input  [31:0] io_RegFileData,
  input  [31:0] io_rsData,
  output [31:0] io_CSROut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] CSReg_0; // @[CSR.scala 23:22]
  reg [31:0] CSReg_1; // @[CSR.scala 23:22]
  reg [31:0] CSReg_2; // @[CSR.scala 23:22]
  reg [31:0] CSReg_3; // @[CSR.scala 23:22]
  reg [31:0] CSReg_4; // @[CSR.scala 23:22]
  reg [31:0] CSReg_5; // @[CSR.scala 23:22]
  reg [31:0] CSReg_6; // @[CSR.scala 23:22]
  reg [31:0] CSReg_7; // @[CSR.scala 23:22]
  reg [31:0] CSReg_8; // @[CSR.scala 23:22]
  reg [31:0] CSReg_9; // @[CSR.scala 23:22]
  reg [31:0] CSReg_10; // @[CSR.scala 23:22]
  reg [31:0] CSReg_11; // @[CSR.scala 23:22]
  reg [31:0] CSReg_12; // @[CSR.scala 23:22]
  reg [31:0] CSReg_13; // @[CSR.scala 23:22]
  reg [31:0] CSReg_14; // @[CSR.scala 23:22]
  reg [31:0] CSReg_15; // @[CSR.scala 23:22]
  reg [31:0] CSReg_16; // @[CSR.scala 23:22]
  reg [31:0] CSReg_17; // @[CSR.scala 23:22]
  reg [31:0] CSReg_18; // @[CSR.scala 23:22]
  reg [31:0] CSReg_19; // @[CSR.scala 23:22]
  reg [31:0] CSReg_20; // @[CSR.scala 23:22]
  reg [31:0] CSReg_21; // @[CSR.scala 23:22]
  reg [31:0] CSReg_22; // @[CSR.scala 23:22]
  reg [31:0] CSReg_23; // @[CSR.scala 23:22]
  reg [31:0] CSReg_24; // @[CSR.scala 23:22]
  reg [31:0] CSReg_25; // @[CSR.scala 23:22]
  reg [31:0] CSReg_26; // @[CSR.scala 23:22]
  reg [31:0] CSReg_27; // @[CSR.scala 23:22]
  reg [31:0] CSReg_28; // @[CSR.scala 23:22]
  reg [31:0] CSReg_29; // @[CSR.scala 23:22]
  reg [31:0] CSReg_30; // @[CSR.scala 23:22]
  reg [31:0] CSReg_31; // @[CSR.scala 23:22]
  reg [31:0] CSReg_32; // @[CSR.scala 23:22]
  reg [31:0] CSReg_33; // @[CSR.scala 23:22]
  reg [31:0] CSReg_34; // @[CSR.scala 23:22]
  reg [31:0] CSReg_35; // @[CSR.scala 23:22]
  reg [31:0] CSReg_36; // @[CSR.scala 23:22]
  reg [31:0] CSReg_37; // @[CSR.scala 23:22]
  reg [31:0] CSReg_38; // @[CSR.scala 23:22]
  reg [31:0] CSReg_39; // @[CSR.scala 23:22]
  reg [31:0] CSReg_40; // @[CSR.scala 23:22]
  reg [31:0] CSReg_41; // @[CSR.scala 23:22]
  reg [31:0] CSReg_42; // @[CSR.scala 23:22]
  reg [31:0] CSReg_43; // @[CSR.scala 23:22]
  reg [31:0] CSReg_44; // @[CSR.scala 23:22]
  reg [31:0] CSReg_45; // @[CSR.scala 23:22]
  reg [31:0] CSReg_46; // @[CSR.scala 23:22]
  reg [31:0] CSReg_47; // @[CSR.scala 23:22]
  reg [31:0] CSReg_48; // @[CSR.scala 23:22]
  reg [31:0] CSReg_49; // @[CSR.scala 23:22]
  reg [31:0] CSReg_50; // @[CSR.scala 23:22]
  reg [31:0] CSReg_51; // @[CSR.scala 23:22]
  reg [31:0] CSReg_52; // @[CSR.scala 23:22]
  reg [31:0] CSReg_53; // @[CSR.scala 23:22]
  reg [31:0] CSReg_54; // @[CSR.scala 23:22]
  reg [31:0] CSReg_55; // @[CSR.scala 23:22]
  reg [31:0] CSReg_56; // @[CSR.scala 23:22]
  reg [31:0] CSReg_57; // @[CSR.scala 23:22]
  reg [31:0] CSReg_58; // @[CSR.scala 23:22]
  reg [31:0] CSReg_59; // @[CSR.scala 23:22]
  reg [31:0] CSReg_60; // @[CSR.scala 23:22]
  reg [31:0] CSReg_61; // @[CSR.scala 23:22]
  reg [31:0] CSReg_62; // @[CSR.scala 23:22]
  reg [31:0] CSReg_63; // @[CSR.scala 23:22]
  reg [31:0] out; // @[CSR.scala 25:20]
  wire [31:0] _GEN_1 = 6'h1 == io_CSRAddr[5:0] ? CSReg_1 : CSReg_0; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_2 = 6'h2 == io_CSRAddr[5:0] ? CSReg_2 : _GEN_1; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_3 = 6'h3 == io_CSRAddr[5:0] ? CSReg_3 : _GEN_2; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_4 = 6'h4 == io_CSRAddr[5:0] ? CSReg_4 : _GEN_3; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_5 = 6'h5 == io_CSRAddr[5:0] ? CSReg_5 : _GEN_4; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_6 = 6'h6 == io_CSRAddr[5:0] ? CSReg_6 : _GEN_5; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_7 = 6'h7 == io_CSRAddr[5:0] ? CSReg_7 : _GEN_6; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_8 = 6'h8 == io_CSRAddr[5:0] ? CSReg_8 : _GEN_7; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_9 = 6'h9 == io_CSRAddr[5:0] ? CSReg_9 : _GEN_8; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_10 = 6'ha == io_CSRAddr[5:0] ? CSReg_10 : _GEN_9; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_11 = 6'hb == io_CSRAddr[5:0] ? CSReg_11 : _GEN_10; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_12 = 6'hc == io_CSRAddr[5:0] ? CSReg_12 : _GEN_11; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_13 = 6'hd == io_CSRAddr[5:0] ? CSReg_13 : _GEN_12; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_14 = 6'he == io_CSRAddr[5:0] ? CSReg_14 : _GEN_13; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_15 = 6'hf == io_CSRAddr[5:0] ? CSReg_15 : _GEN_14; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_16 = 6'h10 == io_CSRAddr[5:0] ? CSReg_16 : _GEN_15; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_17 = 6'h11 == io_CSRAddr[5:0] ? CSReg_17 : _GEN_16; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_18 = 6'h12 == io_CSRAddr[5:0] ? CSReg_18 : _GEN_17; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_19 = 6'h13 == io_CSRAddr[5:0] ? CSReg_19 : _GEN_18; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_20 = 6'h14 == io_CSRAddr[5:0] ? CSReg_20 : _GEN_19; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_21 = 6'h15 == io_CSRAddr[5:0] ? CSReg_21 : _GEN_20; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_22 = 6'h16 == io_CSRAddr[5:0] ? CSReg_22 : _GEN_21; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_23 = 6'h17 == io_CSRAddr[5:0] ? CSReg_23 : _GEN_22; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_24 = 6'h18 == io_CSRAddr[5:0] ? CSReg_24 : _GEN_23; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_25 = 6'h19 == io_CSRAddr[5:0] ? CSReg_25 : _GEN_24; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_26 = 6'h1a == io_CSRAddr[5:0] ? CSReg_26 : _GEN_25; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_27 = 6'h1b == io_CSRAddr[5:0] ? CSReg_27 : _GEN_26; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_28 = 6'h1c == io_CSRAddr[5:0] ? CSReg_28 : _GEN_27; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_29 = 6'h1d == io_CSRAddr[5:0] ? CSReg_29 : _GEN_28; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_30 = 6'h1e == io_CSRAddr[5:0] ? CSReg_30 : _GEN_29; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_31 = 6'h1f == io_CSRAddr[5:0] ? CSReg_31 : _GEN_30; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_32 = 6'h20 == io_CSRAddr[5:0] ? CSReg_32 : _GEN_31; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_33 = 6'h21 == io_CSRAddr[5:0] ? CSReg_33 : _GEN_32; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_34 = 6'h22 == io_CSRAddr[5:0] ? CSReg_34 : _GEN_33; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_35 = 6'h23 == io_CSRAddr[5:0] ? CSReg_35 : _GEN_34; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_36 = 6'h24 == io_CSRAddr[5:0] ? CSReg_36 : _GEN_35; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_37 = 6'h25 == io_CSRAddr[5:0] ? CSReg_37 : _GEN_36; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_38 = 6'h26 == io_CSRAddr[5:0] ? CSReg_38 : _GEN_37; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_39 = 6'h27 == io_CSRAddr[5:0] ? CSReg_39 : _GEN_38; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_40 = 6'h28 == io_CSRAddr[5:0] ? CSReg_40 : _GEN_39; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_41 = 6'h29 == io_CSRAddr[5:0] ? CSReg_41 : _GEN_40; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_42 = 6'h2a == io_CSRAddr[5:0] ? CSReg_42 : _GEN_41; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_43 = 6'h2b == io_CSRAddr[5:0] ? CSReg_43 : _GEN_42; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_44 = 6'h2c == io_CSRAddr[5:0] ? CSReg_44 : _GEN_43; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_45 = 6'h2d == io_CSRAddr[5:0] ? CSReg_45 : _GEN_44; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_46 = 6'h2e == io_CSRAddr[5:0] ? CSReg_46 : _GEN_45; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_47 = 6'h2f == io_CSRAddr[5:0] ? CSReg_47 : _GEN_46; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_48 = 6'h30 == io_CSRAddr[5:0] ? CSReg_48 : _GEN_47; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_49 = 6'h31 == io_CSRAddr[5:0] ? CSReg_49 : _GEN_48; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_50 = 6'h32 == io_CSRAddr[5:0] ? CSReg_50 : _GEN_49; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_51 = 6'h33 == io_CSRAddr[5:0] ? CSReg_51 : _GEN_50; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_52 = 6'h34 == io_CSRAddr[5:0] ? CSReg_52 : _GEN_51; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_53 = 6'h35 == io_CSRAddr[5:0] ? CSReg_53 : _GEN_52; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_54 = 6'h36 == io_CSRAddr[5:0] ? CSReg_54 : _GEN_53; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_55 = 6'h37 == io_CSRAddr[5:0] ? CSReg_55 : _GEN_54; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_56 = 6'h38 == io_CSRAddr[5:0] ? CSReg_56 : _GEN_55; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_57 = 6'h39 == io_CSRAddr[5:0] ? CSReg_57 : _GEN_56; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_58 = 6'h3a == io_CSRAddr[5:0] ? CSReg_58 : _GEN_57; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_59 = 6'h3b == io_CSRAddr[5:0] ? CSReg_59 : _GEN_58; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_60 = 6'h3c == io_CSRAddr[5:0] ? CSReg_60 : _GEN_59; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_61 = 6'h3d == io_CSRAddr[5:0] ? CSReg_61 : _GEN_60; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_62 = 6'h3e == io_CSRAddr[5:0] ? CSReg_62 : _GEN_61; // @[CSR.scala 32:{11,11}]
  wire [31:0] _GEN_63 = 6'h3f == io_CSRAddr[5:0] ? CSReg_63 : _GEN_62; // @[CSR.scala 32:{11,11}]
  wire [31:0] _CSReg_T_1 = _GEN_63 | io_RegFileData; // @[CSR.scala 37:46]
  wire [31:0] _GEN_256 = 6'h0 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_0; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_257 = 6'h1 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_1; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_258 = 6'h2 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_2; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_259 = 6'h3 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_3; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_260 = 6'h4 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_4; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_261 = 6'h5 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_5; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_262 = 6'h6 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_6; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_263 = 6'h7 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_7; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_264 = 6'h8 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_8; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_265 = 6'h9 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_9; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_266 = 6'ha == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_10; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_267 = 6'hb == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_11; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_268 = 6'hc == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_12; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_269 = 6'hd == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_13; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_270 = 6'he == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_14; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_271 = 6'hf == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_15; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_272 = 6'h10 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_16; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_273 = 6'h11 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_17; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_274 = 6'h12 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_18; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_275 = 6'h13 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_19; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_276 = 6'h14 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_20; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_277 = 6'h15 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_21; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_278 = 6'h16 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_22; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_279 = 6'h17 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_23; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_280 = 6'h18 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_24; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_281 = 6'h19 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_25; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_282 = 6'h1a == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_26; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_283 = 6'h1b == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_27; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_284 = 6'h1c == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_28; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_285 = 6'h1d == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_29; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_286 = 6'h1e == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_30; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_287 = 6'h1f == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_31; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_288 = 6'h20 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_32; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_289 = 6'h21 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_33; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_290 = 6'h22 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_34; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_291 = 6'h23 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_35; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_292 = 6'h24 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_36; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_293 = 6'h25 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_37; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_294 = 6'h26 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_38; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_295 = 6'h27 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_39; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_296 = 6'h28 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_40; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_297 = 6'h29 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_41; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_298 = 6'h2a == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_42; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_299 = 6'h2b == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_43; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_300 = 6'h2c == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_44; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_301 = 6'h2d == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_45; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_302 = 6'h2e == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_46; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_303 = 6'h2f == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_47; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_304 = 6'h30 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_48; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_305 = 6'h31 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_49; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_306 = 6'h32 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_50; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_307 = 6'h33 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_51; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_308 = 6'h34 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_52; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_309 = 6'h35 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_53; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_310 = 6'h36 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_54; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_311 = 6'h37 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_55; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_312 = 6'h38 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_56; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_313 = 6'h39 == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_57; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_314 = 6'h3a == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_58; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_315 = 6'h3b == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_59; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_316 = 6'h3c == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_60; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_317 = 6'h3d == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_61; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_318 = 6'h3e == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_62; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _GEN_319 = 6'h3f == io_CSRAddr[5:0] ? _CSReg_T_1 : CSReg_63; // @[CSR.scala 23:22 37:{25,25}]
  wire [31:0] _CSReg_T_3 = ~io_RegFileData; // @[CSR.scala 41:49]
  wire [31:0] _CSReg_T_4 = _GEN_63 & _CSReg_T_3; // @[CSR.scala 41:46]
  wire [31:0] _GEN_448 = 6'h0 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_0; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_449 = 6'h1 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_1; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_450 = 6'h2 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_2; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_451 = 6'h3 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_3; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_452 = 6'h4 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_4; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_453 = 6'h5 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_5; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_454 = 6'h6 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_6; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_455 = 6'h7 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_7; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_456 = 6'h8 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_8; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_457 = 6'h9 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_9; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_458 = 6'ha == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_10; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_459 = 6'hb == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_11; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_460 = 6'hc == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_12; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_461 = 6'hd == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_13; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_462 = 6'he == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_14; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_463 = 6'hf == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_15; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_464 = 6'h10 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_16; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_465 = 6'h11 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_17; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_466 = 6'h12 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_18; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_467 = 6'h13 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_19; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_468 = 6'h14 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_20; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_469 = 6'h15 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_21; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_470 = 6'h16 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_22; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_471 = 6'h17 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_23; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_472 = 6'h18 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_24; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_473 = 6'h19 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_25; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_474 = 6'h1a == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_26; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_475 = 6'h1b == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_27; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_476 = 6'h1c == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_28; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_477 = 6'h1d == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_29; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_478 = 6'h1e == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_30; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_479 = 6'h1f == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_31; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_480 = 6'h20 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_32; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_481 = 6'h21 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_33; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_482 = 6'h22 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_34; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_483 = 6'h23 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_35; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_484 = 6'h24 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_36; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_485 = 6'h25 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_37; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_486 = 6'h26 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_38; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_487 = 6'h27 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_39; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_488 = 6'h28 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_40; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_489 = 6'h29 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_41; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_490 = 6'h2a == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_42; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_491 = 6'h2b == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_43; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_492 = 6'h2c == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_44; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_493 = 6'h2d == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_45; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_494 = 6'h2e == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_46; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_495 = 6'h2f == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_47; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_496 = 6'h30 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_48; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_497 = 6'h31 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_49; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_498 = 6'h32 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_50; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_499 = 6'h33 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_51; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_500 = 6'h34 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_52; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_501 = 6'h35 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_53; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_502 = 6'h36 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_54; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_503 = 6'h37 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_55; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_504 = 6'h38 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_56; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_505 = 6'h39 == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_57; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_506 = 6'h3a == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_58; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_507 = 6'h3b == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_59; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_508 = 6'h3c == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_60; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_509 = 6'h3d == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_61; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_510 = 6'h3e == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_62; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_511 = 6'h3f == io_CSRAddr[5:0] ? _CSReg_T_4 : CSReg_63; // @[CSR.scala 23:22 41:{25,25}]
  wire [31:0] _GEN_576 = 6'h0 == io_CSRAddr[5:0] ? io_rsData : CSReg_0; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_577 = 6'h1 == io_CSRAddr[5:0] ? io_rsData : CSReg_1; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_578 = 6'h2 == io_CSRAddr[5:0] ? io_rsData : CSReg_2; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_579 = 6'h3 == io_CSRAddr[5:0] ? io_rsData : CSReg_3; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_580 = 6'h4 == io_CSRAddr[5:0] ? io_rsData : CSReg_4; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_581 = 6'h5 == io_CSRAddr[5:0] ? io_rsData : CSReg_5; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_582 = 6'h6 == io_CSRAddr[5:0] ? io_rsData : CSReg_6; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_583 = 6'h7 == io_CSRAddr[5:0] ? io_rsData : CSReg_7; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_584 = 6'h8 == io_CSRAddr[5:0] ? io_rsData : CSReg_8; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_585 = 6'h9 == io_CSRAddr[5:0] ? io_rsData : CSReg_9; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_586 = 6'ha == io_CSRAddr[5:0] ? io_rsData : CSReg_10; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_587 = 6'hb == io_CSRAddr[5:0] ? io_rsData : CSReg_11; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_588 = 6'hc == io_CSRAddr[5:0] ? io_rsData : CSReg_12; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_589 = 6'hd == io_CSRAddr[5:0] ? io_rsData : CSReg_13; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_590 = 6'he == io_CSRAddr[5:0] ? io_rsData : CSReg_14; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_591 = 6'hf == io_CSRAddr[5:0] ? io_rsData : CSReg_15; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_592 = 6'h10 == io_CSRAddr[5:0] ? io_rsData : CSReg_16; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_593 = 6'h11 == io_CSRAddr[5:0] ? io_rsData : CSReg_17; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_594 = 6'h12 == io_CSRAddr[5:0] ? io_rsData : CSReg_18; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_595 = 6'h13 == io_CSRAddr[5:0] ? io_rsData : CSReg_19; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_596 = 6'h14 == io_CSRAddr[5:0] ? io_rsData : CSReg_20; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_597 = 6'h15 == io_CSRAddr[5:0] ? io_rsData : CSReg_21; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_598 = 6'h16 == io_CSRAddr[5:0] ? io_rsData : CSReg_22; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_599 = 6'h17 == io_CSRAddr[5:0] ? io_rsData : CSReg_23; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_600 = 6'h18 == io_CSRAddr[5:0] ? io_rsData : CSReg_24; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_601 = 6'h19 == io_CSRAddr[5:0] ? io_rsData : CSReg_25; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_602 = 6'h1a == io_CSRAddr[5:0] ? io_rsData : CSReg_26; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_603 = 6'h1b == io_CSRAddr[5:0] ? io_rsData : CSReg_27; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_604 = 6'h1c == io_CSRAddr[5:0] ? io_rsData : CSReg_28; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_605 = 6'h1d == io_CSRAddr[5:0] ? io_rsData : CSReg_29; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_606 = 6'h1e == io_CSRAddr[5:0] ? io_rsData : CSReg_30; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_607 = 6'h1f == io_CSRAddr[5:0] ? io_rsData : CSReg_31; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_608 = 6'h20 == io_CSRAddr[5:0] ? io_rsData : CSReg_32; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_609 = 6'h21 == io_CSRAddr[5:0] ? io_rsData : CSReg_33; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_610 = 6'h22 == io_CSRAddr[5:0] ? io_rsData : CSReg_34; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_611 = 6'h23 == io_CSRAddr[5:0] ? io_rsData : CSReg_35; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_612 = 6'h24 == io_CSRAddr[5:0] ? io_rsData : CSReg_36; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_613 = 6'h25 == io_CSRAddr[5:0] ? io_rsData : CSReg_37; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_614 = 6'h26 == io_CSRAddr[5:0] ? io_rsData : CSReg_38; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_615 = 6'h27 == io_CSRAddr[5:0] ? io_rsData : CSReg_39; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_616 = 6'h28 == io_CSRAddr[5:0] ? io_rsData : CSReg_40; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_617 = 6'h29 == io_CSRAddr[5:0] ? io_rsData : CSReg_41; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_618 = 6'h2a == io_CSRAddr[5:0] ? io_rsData : CSReg_42; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_619 = 6'h2b == io_CSRAddr[5:0] ? io_rsData : CSReg_43; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_620 = 6'h2c == io_CSRAddr[5:0] ? io_rsData : CSReg_44; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_621 = 6'h2d == io_CSRAddr[5:0] ? io_rsData : CSReg_45; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_622 = 6'h2e == io_CSRAddr[5:0] ? io_rsData : CSReg_46; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_623 = 6'h2f == io_CSRAddr[5:0] ? io_rsData : CSReg_47; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_624 = 6'h30 == io_CSRAddr[5:0] ? io_rsData : CSReg_48; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_625 = 6'h31 == io_CSRAddr[5:0] ? io_rsData : CSReg_49; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_626 = 6'h32 == io_CSRAddr[5:0] ? io_rsData : CSReg_50; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_627 = 6'h33 == io_CSRAddr[5:0] ? io_rsData : CSReg_51; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_628 = 6'h34 == io_CSRAddr[5:0] ? io_rsData : CSReg_52; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_629 = 6'h35 == io_CSRAddr[5:0] ? io_rsData : CSReg_53; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_630 = 6'h36 == io_CSRAddr[5:0] ? io_rsData : CSReg_54; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_631 = 6'h37 == io_CSRAddr[5:0] ? io_rsData : CSReg_55; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_632 = 6'h38 == io_CSRAddr[5:0] ? io_rsData : CSReg_56; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_633 = 6'h39 == io_CSRAddr[5:0] ? io_rsData : CSReg_57; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_634 = 6'h3a == io_CSRAddr[5:0] ? io_rsData : CSReg_58; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_635 = 6'h3b == io_CSRAddr[5:0] ? io_rsData : CSReg_59; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_636 = 6'h3c == io_CSRAddr[5:0] ? io_rsData : CSReg_60; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_637 = 6'h3d == io_CSRAddr[5:0] ? io_rsData : CSReg_61; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_638 = 6'h3e == io_CSRAddr[5:0] ? io_rsData : CSReg_62; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _GEN_639 = 6'h3f == io_CSRAddr[5:0] ? io_rsData : CSReg_63; // @[CSR.scala 23:22 45:{25,25}]
  wire [31:0] _CSReg_T_6 = _GEN_63 | io_rsData; // @[CSR.scala 49:46]
  wire [31:0] _GEN_768 = 6'h0 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_0; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_769 = 6'h1 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_1; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_770 = 6'h2 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_2; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_771 = 6'h3 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_3; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_772 = 6'h4 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_4; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_773 = 6'h5 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_5; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_774 = 6'h6 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_6; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_775 = 6'h7 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_7; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_776 = 6'h8 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_8; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_777 = 6'h9 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_9; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_778 = 6'ha == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_10; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_779 = 6'hb == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_11; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_780 = 6'hc == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_12; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_781 = 6'hd == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_13; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_782 = 6'he == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_14; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_783 = 6'hf == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_15; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_784 = 6'h10 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_16; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_785 = 6'h11 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_17; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_786 = 6'h12 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_18; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_787 = 6'h13 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_19; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_788 = 6'h14 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_20; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_789 = 6'h15 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_21; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_790 = 6'h16 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_22; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_791 = 6'h17 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_23; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_792 = 6'h18 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_24; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_793 = 6'h19 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_25; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_794 = 6'h1a == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_26; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_795 = 6'h1b == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_27; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_796 = 6'h1c == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_28; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_797 = 6'h1d == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_29; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_798 = 6'h1e == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_30; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_799 = 6'h1f == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_31; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_800 = 6'h20 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_32; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_801 = 6'h21 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_33; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_802 = 6'h22 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_34; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_803 = 6'h23 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_35; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_804 = 6'h24 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_36; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_805 = 6'h25 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_37; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_806 = 6'h26 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_38; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_807 = 6'h27 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_39; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_808 = 6'h28 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_40; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_809 = 6'h29 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_41; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_810 = 6'h2a == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_42; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_811 = 6'h2b == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_43; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_812 = 6'h2c == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_44; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_813 = 6'h2d == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_45; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_814 = 6'h2e == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_46; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_815 = 6'h2f == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_47; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_816 = 6'h30 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_48; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_817 = 6'h31 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_49; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_818 = 6'h32 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_50; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_819 = 6'h33 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_51; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_820 = 6'h34 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_52; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_821 = 6'h35 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_53; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_822 = 6'h36 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_54; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_823 = 6'h37 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_55; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_824 = 6'h38 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_56; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_825 = 6'h39 == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_57; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_826 = 6'h3a == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_58; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_827 = 6'h3b == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_59; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_828 = 6'h3c == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_60; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_829 = 6'h3d == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_61; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_830 = 6'h3e == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_62; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _GEN_831 = 6'h3f == io_CSRAddr[5:0] ? _CSReg_T_6 : CSReg_63; // @[CSR.scala 23:22 49:{25,25}]
  wire [31:0] _CSReg_T_8 = ~io_rsData; // @[CSR.scala 53:49]
  wire [31:0] _CSReg_T_9 = _GEN_63 & _CSReg_T_8; // @[CSR.scala 53:46]
  wire [31:0] _GEN_960 = 6'h0 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_0; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_961 = 6'h1 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_1; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_962 = 6'h2 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_2; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_963 = 6'h3 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_3; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_964 = 6'h4 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_4; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_965 = 6'h5 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_5; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_966 = 6'h6 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_6; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_967 = 6'h7 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_7; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_968 = 6'h8 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_8; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_969 = 6'h9 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_9; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_970 = 6'ha == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_10; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_971 = 6'hb == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_11; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_972 = 6'hc == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_12; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_973 = 6'hd == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_13; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_974 = 6'he == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_14; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_975 = 6'hf == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_15; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_976 = 6'h10 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_16; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_977 = 6'h11 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_17; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_978 = 6'h12 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_18; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_979 = 6'h13 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_19; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_980 = 6'h14 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_20; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_981 = 6'h15 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_21; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_982 = 6'h16 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_22; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_983 = 6'h17 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_23; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_984 = 6'h18 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_24; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_985 = 6'h19 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_25; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_986 = 6'h1a == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_26; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_987 = 6'h1b == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_27; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_988 = 6'h1c == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_28; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_989 = 6'h1d == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_29; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_990 = 6'h1e == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_30; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_991 = 6'h1f == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_31; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_992 = 6'h20 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_32; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_993 = 6'h21 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_33; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_994 = 6'h22 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_34; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_995 = 6'h23 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_35; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_996 = 6'h24 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_36; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_997 = 6'h25 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_37; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_998 = 6'h26 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_38; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_999 = 6'h27 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_39; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1000 = 6'h28 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_40; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1001 = 6'h29 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_41; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1002 = 6'h2a == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_42; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1003 = 6'h2b == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_43; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1004 = 6'h2c == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_44; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1005 = 6'h2d == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_45; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1006 = 6'h2e == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_46; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1007 = 6'h2f == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_47; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1008 = 6'h30 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_48; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1009 = 6'h31 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_49; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1010 = 6'h32 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_50; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1011 = 6'h33 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_51; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1012 = 6'h34 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_52; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1013 = 6'h35 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_53; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1014 = 6'h36 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_54; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1015 = 6'h37 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_55; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1016 = 6'h38 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_56; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1017 = 6'h39 == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_57; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1018 = 6'h3a == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_58; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1019 = 6'h3b == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_59; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1020 = 6'h3c == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_60; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1021 = 6'h3d == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_61; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1022 = 6'h3e == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_62; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1023 = 6'h3f == io_CSRAddr[5:0] ? _CSReg_T_9 : CSReg_63; // @[CSR.scala 23:22 53:{25,25}]
  wire [31:0] _GEN_1024 = 3'h6 == io_CSRType ? _GEN_63 : out; // @[CSR.scala 27:21 52:11 25:20]
  wire [31:0] _GEN_1025 = 3'h6 == io_CSRType ? _GEN_960 : CSReg_0; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1026 = 3'h6 == io_CSRType ? _GEN_961 : CSReg_1; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1027 = 3'h6 == io_CSRType ? _GEN_962 : CSReg_2; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1028 = 3'h6 == io_CSRType ? _GEN_963 : CSReg_3; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1029 = 3'h6 == io_CSRType ? _GEN_964 : CSReg_4; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1030 = 3'h6 == io_CSRType ? _GEN_965 : CSReg_5; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1031 = 3'h6 == io_CSRType ? _GEN_966 : CSReg_6; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1032 = 3'h6 == io_CSRType ? _GEN_967 : CSReg_7; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1033 = 3'h6 == io_CSRType ? _GEN_968 : CSReg_8; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1034 = 3'h6 == io_CSRType ? _GEN_969 : CSReg_9; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1035 = 3'h6 == io_CSRType ? _GEN_970 : CSReg_10; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1036 = 3'h6 == io_CSRType ? _GEN_971 : CSReg_11; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1037 = 3'h6 == io_CSRType ? _GEN_972 : CSReg_12; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1038 = 3'h6 == io_CSRType ? _GEN_973 : CSReg_13; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1039 = 3'h6 == io_CSRType ? _GEN_974 : CSReg_14; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1040 = 3'h6 == io_CSRType ? _GEN_975 : CSReg_15; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1041 = 3'h6 == io_CSRType ? _GEN_976 : CSReg_16; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1042 = 3'h6 == io_CSRType ? _GEN_977 : CSReg_17; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1043 = 3'h6 == io_CSRType ? _GEN_978 : CSReg_18; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1044 = 3'h6 == io_CSRType ? _GEN_979 : CSReg_19; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1045 = 3'h6 == io_CSRType ? _GEN_980 : CSReg_20; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1046 = 3'h6 == io_CSRType ? _GEN_981 : CSReg_21; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1047 = 3'h6 == io_CSRType ? _GEN_982 : CSReg_22; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1048 = 3'h6 == io_CSRType ? _GEN_983 : CSReg_23; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1049 = 3'h6 == io_CSRType ? _GEN_984 : CSReg_24; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1050 = 3'h6 == io_CSRType ? _GEN_985 : CSReg_25; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1051 = 3'h6 == io_CSRType ? _GEN_986 : CSReg_26; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1052 = 3'h6 == io_CSRType ? _GEN_987 : CSReg_27; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1053 = 3'h6 == io_CSRType ? _GEN_988 : CSReg_28; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1054 = 3'h6 == io_CSRType ? _GEN_989 : CSReg_29; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1055 = 3'h6 == io_CSRType ? _GEN_990 : CSReg_30; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1056 = 3'h6 == io_CSRType ? _GEN_991 : CSReg_31; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1057 = 3'h6 == io_CSRType ? _GEN_992 : CSReg_32; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1058 = 3'h6 == io_CSRType ? _GEN_993 : CSReg_33; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1059 = 3'h6 == io_CSRType ? _GEN_994 : CSReg_34; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1060 = 3'h6 == io_CSRType ? _GEN_995 : CSReg_35; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1061 = 3'h6 == io_CSRType ? _GEN_996 : CSReg_36; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1062 = 3'h6 == io_CSRType ? _GEN_997 : CSReg_37; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1063 = 3'h6 == io_CSRType ? _GEN_998 : CSReg_38; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1064 = 3'h6 == io_CSRType ? _GEN_999 : CSReg_39; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1065 = 3'h6 == io_CSRType ? _GEN_1000 : CSReg_40; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1066 = 3'h6 == io_CSRType ? _GEN_1001 : CSReg_41; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1067 = 3'h6 == io_CSRType ? _GEN_1002 : CSReg_42; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1068 = 3'h6 == io_CSRType ? _GEN_1003 : CSReg_43; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1069 = 3'h6 == io_CSRType ? _GEN_1004 : CSReg_44; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1070 = 3'h6 == io_CSRType ? _GEN_1005 : CSReg_45; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1071 = 3'h6 == io_CSRType ? _GEN_1006 : CSReg_46; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1072 = 3'h6 == io_CSRType ? _GEN_1007 : CSReg_47; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1073 = 3'h6 == io_CSRType ? _GEN_1008 : CSReg_48; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1074 = 3'h6 == io_CSRType ? _GEN_1009 : CSReg_49; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1075 = 3'h6 == io_CSRType ? _GEN_1010 : CSReg_50; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1076 = 3'h6 == io_CSRType ? _GEN_1011 : CSReg_51; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1077 = 3'h6 == io_CSRType ? _GEN_1012 : CSReg_52; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1078 = 3'h6 == io_CSRType ? _GEN_1013 : CSReg_53; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1079 = 3'h6 == io_CSRType ? _GEN_1014 : CSReg_54; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1080 = 3'h6 == io_CSRType ? _GEN_1015 : CSReg_55; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1081 = 3'h6 == io_CSRType ? _GEN_1016 : CSReg_56; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1082 = 3'h6 == io_CSRType ? _GEN_1017 : CSReg_57; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1083 = 3'h6 == io_CSRType ? _GEN_1018 : CSReg_58; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1084 = 3'h6 == io_CSRType ? _GEN_1019 : CSReg_59; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1085 = 3'h6 == io_CSRType ? _GEN_1020 : CSReg_60; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1086 = 3'h6 == io_CSRType ? _GEN_1021 : CSReg_61; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1087 = 3'h6 == io_CSRType ? _GEN_1022 : CSReg_62; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1088 = 3'h6 == io_CSRType ? _GEN_1023 : CSReg_63; // @[CSR.scala 27:21 23:22]
  wire [31:0] _GEN_1089 = 3'h5 == io_CSRType ? _GEN_63 : _GEN_1024; // @[CSR.scala 27:21 48:11]
  wire [31:0] _GEN_1090 = 3'h5 == io_CSRType ? _GEN_768 : _GEN_1025; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1091 = 3'h5 == io_CSRType ? _GEN_769 : _GEN_1026; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1092 = 3'h5 == io_CSRType ? _GEN_770 : _GEN_1027; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1093 = 3'h5 == io_CSRType ? _GEN_771 : _GEN_1028; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1094 = 3'h5 == io_CSRType ? _GEN_772 : _GEN_1029; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1095 = 3'h5 == io_CSRType ? _GEN_773 : _GEN_1030; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1096 = 3'h5 == io_CSRType ? _GEN_774 : _GEN_1031; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1097 = 3'h5 == io_CSRType ? _GEN_775 : _GEN_1032; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1098 = 3'h5 == io_CSRType ? _GEN_776 : _GEN_1033; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1099 = 3'h5 == io_CSRType ? _GEN_777 : _GEN_1034; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1100 = 3'h5 == io_CSRType ? _GEN_778 : _GEN_1035; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1101 = 3'h5 == io_CSRType ? _GEN_779 : _GEN_1036; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1102 = 3'h5 == io_CSRType ? _GEN_780 : _GEN_1037; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1103 = 3'h5 == io_CSRType ? _GEN_781 : _GEN_1038; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1104 = 3'h5 == io_CSRType ? _GEN_782 : _GEN_1039; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1105 = 3'h5 == io_CSRType ? _GEN_783 : _GEN_1040; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1106 = 3'h5 == io_CSRType ? _GEN_784 : _GEN_1041; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1107 = 3'h5 == io_CSRType ? _GEN_785 : _GEN_1042; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1108 = 3'h5 == io_CSRType ? _GEN_786 : _GEN_1043; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1109 = 3'h5 == io_CSRType ? _GEN_787 : _GEN_1044; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1110 = 3'h5 == io_CSRType ? _GEN_788 : _GEN_1045; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1111 = 3'h5 == io_CSRType ? _GEN_789 : _GEN_1046; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1112 = 3'h5 == io_CSRType ? _GEN_790 : _GEN_1047; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1113 = 3'h5 == io_CSRType ? _GEN_791 : _GEN_1048; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1114 = 3'h5 == io_CSRType ? _GEN_792 : _GEN_1049; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1115 = 3'h5 == io_CSRType ? _GEN_793 : _GEN_1050; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1116 = 3'h5 == io_CSRType ? _GEN_794 : _GEN_1051; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1117 = 3'h5 == io_CSRType ? _GEN_795 : _GEN_1052; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1118 = 3'h5 == io_CSRType ? _GEN_796 : _GEN_1053; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1119 = 3'h5 == io_CSRType ? _GEN_797 : _GEN_1054; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1120 = 3'h5 == io_CSRType ? _GEN_798 : _GEN_1055; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1121 = 3'h5 == io_CSRType ? _GEN_799 : _GEN_1056; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1122 = 3'h5 == io_CSRType ? _GEN_800 : _GEN_1057; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1123 = 3'h5 == io_CSRType ? _GEN_801 : _GEN_1058; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1124 = 3'h5 == io_CSRType ? _GEN_802 : _GEN_1059; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1125 = 3'h5 == io_CSRType ? _GEN_803 : _GEN_1060; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1126 = 3'h5 == io_CSRType ? _GEN_804 : _GEN_1061; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1127 = 3'h5 == io_CSRType ? _GEN_805 : _GEN_1062; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1128 = 3'h5 == io_CSRType ? _GEN_806 : _GEN_1063; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1129 = 3'h5 == io_CSRType ? _GEN_807 : _GEN_1064; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1130 = 3'h5 == io_CSRType ? _GEN_808 : _GEN_1065; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1131 = 3'h5 == io_CSRType ? _GEN_809 : _GEN_1066; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1132 = 3'h5 == io_CSRType ? _GEN_810 : _GEN_1067; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1133 = 3'h5 == io_CSRType ? _GEN_811 : _GEN_1068; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1134 = 3'h5 == io_CSRType ? _GEN_812 : _GEN_1069; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1135 = 3'h5 == io_CSRType ? _GEN_813 : _GEN_1070; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1136 = 3'h5 == io_CSRType ? _GEN_814 : _GEN_1071; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1137 = 3'h5 == io_CSRType ? _GEN_815 : _GEN_1072; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1138 = 3'h5 == io_CSRType ? _GEN_816 : _GEN_1073; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1139 = 3'h5 == io_CSRType ? _GEN_817 : _GEN_1074; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1140 = 3'h5 == io_CSRType ? _GEN_818 : _GEN_1075; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1141 = 3'h5 == io_CSRType ? _GEN_819 : _GEN_1076; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1142 = 3'h5 == io_CSRType ? _GEN_820 : _GEN_1077; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1143 = 3'h5 == io_CSRType ? _GEN_821 : _GEN_1078; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1144 = 3'h5 == io_CSRType ? _GEN_822 : _GEN_1079; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1145 = 3'h5 == io_CSRType ? _GEN_823 : _GEN_1080; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1146 = 3'h5 == io_CSRType ? _GEN_824 : _GEN_1081; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1147 = 3'h5 == io_CSRType ? _GEN_825 : _GEN_1082; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1148 = 3'h5 == io_CSRType ? _GEN_826 : _GEN_1083; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1149 = 3'h5 == io_CSRType ? _GEN_827 : _GEN_1084; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1150 = 3'h5 == io_CSRType ? _GEN_828 : _GEN_1085; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1151 = 3'h5 == io_CSRType ? _GEN_829 : _GEN_1086; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1152 = 3'h5 == io_CSRType ? _GEN_830 : _GEN_1087; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1153 = 3'h5 == io_CSRType ? _GEN_831 : _GEN_1088; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1154 = 3'h4 == io_CSRType ? _GEN_63 : _GEN_1089; // @[CSR.scala 27:21 44:11]
  wire [31:0] _GEN_1155 = 3'h4 == io_CSRType ? _GEN_576 : _GEN_1090; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1156 = 3'h4 == io_CSRType ? _GEN_577 : _GEN_1091; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1157 = 3'h4 == io_CSRType ? _GEN_578 : _GEN_1092; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1158 = 3'h4 == io_CSRType ? _GEN_579 : _GEN_1093; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1159 = 3'h4 == io_CSRType ? _GEN_580 : _GEN_1094; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1160 = 3'h4 == io_CSRType ? _GEN_581 : _GEN_1095; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1161 = 3'h4 == io_CSRType ? _GEN_582 : _GEN_1096; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1162 = 3'h4 == io_CSRType ? _GEN_583 : _GEN_1097; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1163 = 3'h4 == io_CSRType ? _GEN_584 : _GEN_1098; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1164 = 3'h4 == io_CSRType ? _GEN_585 : _GEN_1099; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1165 = 3'h4 == io_CSRType ? _GEN_586 : _GEN_1100; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1166 = 3'h4 == io_CSRType ? _GEN_587 : _GEN_1101; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1167 = 3'h4 == io_CSRType ? _GEN_588 : _GEN_1102; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1168 = 3'h4 == io_CSRType ? _GEN_589 : _GEN_1103; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1169 = 3'h4 == io_CSRType ? _GEN_590 : _GEN_1104; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1170 = 3'h4 == io_CSRType ? _GEN_591 : _GEN_1105; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1171 = 3'h4 == io_CSRType ? _GEN_592 : _GEN_1106; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1172 = 3'h4 == io_CSRType ? _GEN_593 : _GEN_1107; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1173 = 3'h4 == io_CSRType ? _GEN_594 : _GEN_1108; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1174 = 3'h4 == io_CSRType ? _GEN_595 : _GEN_1109; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1175 = 3'h4 == io_CSRType ? _GEN_596 : _GEN_1110; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1176 = 3'h4 == io_CSRType ? _GEN_597 : _GEN_1111; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1177 = 3'h4 == io_CSRType ? _GEN_598 : _GEN_1112; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1178 = 3'h4 == io_CSRType ? _GEN_599 : _GEN_1113; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1179 = 3'h4 == io_CSRType ? _GEN_600 : _GEN_1114; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1180 = 3'h4 == io_CSRType ? _GEN_601 : _GEN_1115; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1181 = 3'h4 == io_CSRType ? _GEN_602 : _GEN_1116; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1182 = 3'h4 == io_CSRType ? _GEN_603 : _GEN_1117; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1183 = 3'h4 == io_CSRType ? _GEN_604 : _GEN_1118; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1184 = 3'h4 == io_CSRType ? _GEN_605 : _GEN_1119; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1185 = 3'h4 == io_CSRType ? _GEN_606 : _GEN_1120; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1186 = 3'h4 == io_CSRType ? _GEN_607 : _GEN_1121; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1187 = 3'h4 == io_CSRType ? _GEN_608 : _GEN_1122; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1188 = 3'h4 == io_CSRType ? _GEN_609 : _GEN_1123; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1189 = 3'h4 == io_CSRType ? _GEN_610 : _GEN_1124; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1190 = 3'h4 == io_CSRType ? _GEN_611 : _GEN_1125; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1191 = 3'h4 == io_CSRType ? _GEN_612 : _GEN_1126; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1192 = 3'h4 == io_CSRType ? _GEN_613 : _GEN_1127; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1193 = 3'h4 == io_CSRType ? _GEN_614 : _GEN_1128; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1194 = 3'h4 == io_CSRType ? _GEN_615 : _GEN_1129; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1195 = 3'h4 == io_CSRType ? _GEN_616 : _GEN_1130; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1196 = 3'h4 == io_CSRType ? _GEN_617 : _GEN_1131; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1197 = 3'h4 == io_CSRType ? _GEN_618 : _GEN_1132; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1198 = 3'h4 == io_CSRType ? _GEN_619 : _GEN_1133; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1199 = 3'h4 == io_CSRType ? _GEN_620 : _GEN_1134; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1200 = 3'h4 == io_CSRType ? _GEN_621 : _GEN_1135; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1201 = 3'h4 == io_CSRType ? _GEN_622 : _GEN_1136; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1202 = 3'h4 == io_CSRType ? _GEN_623 : _GEN_1137; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1203 = 3'h4 == io_CSRType ? _GEN_624 : _GEN_1138; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1204 = 3'h4 == io_CSRType ? _GEN_625 : _GEN_1139; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1205 = 3'h4 == io_CSRType ? _GEN_626 : _GEN_1140; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1206 = 3'h4 == io_CSRType ? _GEN_627 : _GEN_1141; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1207 = 3'h4 == io_CSRType ? _GEN_628 : _GEN_1142; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1208 = 3'h4 == io_CSRType ? _GEN_629 : _GEN_1143; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1209 = 3'h4 == io_CSRType ? _GEN_630 : _GEN_1144; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1210 = 3'h4 == io_CSRType ? _GEN_631 : _GEN_1145; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1211 = 3'h4 == io_CSRType ? _GEN_632 : _GEN_1146; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1212 = 3'h4 == io_CSRType ? _GEN_633 : _GEN_1147; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1213 = 3'h4 == io_CSRType ? _GEN_634 : _GEN_1148; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1214 = 3'h4 == io_CSRType ? _GEN_635 : _GEN_1149; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1215 = 3'h4 == io_CSRType ? _GEN_636 : _GEN_1150; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1216 = 3'h4 == io_CSRType ? _GEN_637 : _GEN_1151; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1217 = 3'h4 == io_CSRType ? _GEN_638 : _GEN_1152; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1218 = 3'h4 == io_CSRType ? _GEN_639 : _GEN_1153; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1219 = 3'h3 == io_CSRType ? _GEN_63 : _GEN_1154; // @[CSR.scala 27:21 40:11]
  wire [31:0] _GEN_1220 = 3'h3 == io_CSRType ? _GEN_448 : _GEN_1155; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1221 = 3'h3 == io_CSRType ? _GEN_449 : _GEN_1156; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1222 = 3'h3 == io_CSRType ? _GEN_450 : _GEN_1157; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1223 = 3'h3 == io_CSRType ? _GEN_451 : _GEN_1158; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1224 = 3'h3 == io_CSRType ? _GEN_452 : _GEN_1159; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1225 = 3'h3 == io_CSRType ? _GEN_453 : _GEN_1160; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1226 = 3'h3 == io_CSRType ? _GEN_454 : _GEN_1161; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1227 = 3'h3 == io_CSRType ? _GEN_455 : _GEN_1162; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1228 = 3'h3 == io_CSRType ? _GEN_456 : _GEN_1163; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1229 = 3'h3 == io_CSRType ? _GEN_457 : _GEN_1164; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1230 = 3'h3 == io_CSRType ? _GEN_458 : _GEN_1165; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1231 = 3'h3 == io_CSRType ? _GEN_459 : _GEN_1166; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1232 = 3'h3 == io_CSRType ? _GEN_460 : _GEN_1167; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1233 = 3'h3 == io_CSRType ? _GEN_461 : _GEN_1168; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1234 = 3'h3 == io_CSRType ? _GEN_462 : _GEN_1169; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1235 = 3'h3 == io_CSRType ? _GEN_463 : _GEN_1170; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1236 = 3'h3 == io_CSRType ? _GEN_464 : _GEN_1171; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1237 = 3'h3 == io_CSRType ? _GEN_465 : _GEN_1172; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1238 = 3'h3 == io_CSRType ? _GEN_466 : _GEN_1173; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1239 = 3'h3 == io_CSRType ? _GEN_467 : _GEN_1174; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1240 = 3'h3 == io_CSRType ? _GEN_468 : _GEN_1175; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1241 = 3'h3 == io_CSRType ? _GEN_469 : _GEN_1176; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1242 = 3'h3 == io_CSRType ? _GEN_470 : _GEN_1177; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1243 = 3'h3 == io_CSRType ? _GEN_471 : _GEN_1178; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1244 = 3'h3 == io_CSRType ? _GEN_472 : _GEN_1179; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1245 = 3'h3 == io_CSRType ? _GEN_473 : _GEN_1180; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1246 = 3'h3 == io_CSRType ? _GEN_474 : _GEN_1181; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1247 = 3'h3 == io_CSRType ? _GEN_475 : _GEN_1182; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1248 = 3'h3 == io_CSRType ? _GEN_476 : _GEN_1183; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1249 = 3'h3 == io_CSRType ? _GEN_477 : _GEN_1184; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1250 = 3'h3 == io_CSRType ? _GEN_478 : _GEN_1185; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1251 = 3'h3 == io_CSRType ? _GEN_479 : _GEN_1186; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1252 = 3'h3 == io_CSRType ? _GEN_480 : _GEN_1187; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1253 = 3'h3 == io_CSRType ? _GEN_481 : _GEN_1188; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1254 = 3'h3 == io_CSRType ? _GEN_482 : _GEN_1189; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1255 = 3'h3 == io_CSRType ? _GEN_483 : _GEN_1190; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1256 = 3'h3 == io_CSRType ? _GEN_484 : _GEN_1191; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1257 = 3'h3 == io_CSRType ? _GEN_485 : _GEN_1192; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1258 = 3'h3 == io_CSRType ? _GEN_486 : _GEN_1193; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1259 = 3'h3 == io_CSRType ? _GEN_487 : _GEN_1194; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1260 = 3'h3 == io_CSRType ? _GEN_488 : _GEN_1195; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1261 = 3'h3 == io_CSRType ? _GEN_489 : _GEN_1196; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1262 = 3'h3 == io_CSRType ? _GEN_490 : _GEN_1197; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1263 = 3'h3 == io_CSRType ? _GEN_491 : _GEN_1198; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1264 = 3'h3 == io_CSRType ? _GEN_492 : _GEN_1199; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1265 = 3'h3 == io_CSRType ? _GEN_493 : _GEN_1200; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1266 = 3'h3 == io_CSRType ? _GEN_494 : _GEN_1201; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1267 = 3'h3 == io_CSRType ? _GEN_495 : _GEN_1202; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1268 = 3'h3 == io_CSRType ? _GEN_496 : _GEN_1203; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1269 = 3'h3 == io_CSRType ? _GEN_497 : _GEN_1204; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1270 = 3'h3 == io_CSRType ? _GEN_498 : _GEN_1205; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1271 = 3'h3 == io_CSRType ? _GEN_499 : _GEN_1206; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1272 = 3'h3 == io_CSRType ? _GEN_500 : _GEN_1207; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1273 = 3'h3 == io_CSRType ? _GEN_501 : _GEN_1208; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1274 = 3'h3 == io_CSRType ? _GEN_502 : _GEN_1209; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1275 = 3'h3 == io_CSRType ? _GEN_503 : _GEN_1210; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1276 = 3'h3 == io_CSRType ? _GEN_504 : _GEN_1211; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1277 = 3'h3 == io_CSRType ? _GEN_505 : _GEN_1212; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1278 = 3'h3 == io_CSRType ? _GEN_506 : _GEN_1213; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1279 = 3'h3 == io_CSRType ? _GEN_507 : _GEN_1214; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1280 = 3'h3 == io_CSRType ? _GEN_508 : _GEN_1215; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1281 = 3'h3 == io_CSRType ? _GEN_509 : _GEN_1216; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1282 = 3'h3 == io_CSRType ? _GEN_510 : _GEN_1217; // @[CSR.scala 27:21]
  wire [31:0] _GEN_1283 = 3'h3 == io_CSRType ? _GEN_511 : _GEN_1218; // @[CSR.scala 27:21]
  assign io_CSROut = out; // @[CSR.scala 59:13]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_0 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h0 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_0 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_0 <= _GEN_256;
      end else begin
        CSReg_0 <= _GEN_1220;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_1 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_1 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_1 <= _GEN_257;
      end else begin
        CSReg_1 <= _GEN_1221;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_2 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_2 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_2 <= _GEN_258;
      end else begin
        CSReg_2 <= _GEN_1222;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_3 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_3 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_3 <= _GEN_259;
      end else begin
        CSReg_3 <= _GEN_1223;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_4 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h4 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_4 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_4 <= _GEN_260;
      end else begin
        CSReg_4 <= _GEN_1224;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_5 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h5 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_5 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_5 <= _GEN_261;
      end else begin
        CSReg_5 <= _GEN_1225;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_6 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h6 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_6 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_6 <= _GEN_262;
      end else begin
        CSReg_6 <= _GEN_1226;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_7 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h7 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_7 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_7 <= _GEN_263;
      end else begin
        CSReg_7 <= _GEN_1227;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_8 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h8 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_8 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_8 <= _GEN_264;
      end else begin
        CSReg_8 <= _GEN_1228;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_9 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h9 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_9 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_9 <= _GEN_265;
      end else begin
        CSReg_9 <= _GEN_1229;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_10 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'ha == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_10 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_10 <= _GEN_266;
      end else begin
        CSReg_10 <= _GEN_1230;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_11 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'hb == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_11 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_11 <= _GEN_267;
      end else begin
        CSReg_11 <= _GEN_1231;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_12 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'hc == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_12 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_12 <= _GEN_268;
      end else begin
        CSReg_12 <= _GEN_1232;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_13 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'hd == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_13 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_13 <= _GEN_269;
      end else begin
        CSReg_13 <= _GEN_1233;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_14 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'he == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_14 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_14 <= _GEN_270;
      end else begin
        CSReg_14 <= _GEN_1234;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_15 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'hf == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_15 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_15 <= _GEN_271;
      end else begin
        CSReg_15 <= _GEN_1235;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_16 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h10 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_16 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_16 <= _GEN_272;
      end else begin
        CSReg_16 <= _GEN_1236;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_17 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h11 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_17 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_17 <= _GEN_273;
      end else begin
        CSReg_17 <= _GEN_1237;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_18 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h12 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_18 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_18 <= _GEN_274;
      end else begin
        CSReg_18 <= _GEN_1238;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_19 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h13 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_19 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_19 <= _GEN_275;
      end else begin
        CSReg_19 <= _GEN_1239;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_20 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h14 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_20 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_20 <= _GEN_276;
      end else begin
        CSReg_20 <= _GEN_1240;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_21 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h15 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_21 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_21 <= _GEN_277;
      end else begin
        CSReg_21 <= _GEN_1241;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_22 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h16 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_22 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_22 <= _GEN_278;
      end else begin
        CSReg_22 <= _GEN_1242;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_23 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h17 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_23 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_23 <= _GEN_279;
      end else begin
        CSReg_23 <= _GEN_1243;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_24 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h18 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_24 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_24 <= _GEN_280;
      end else begin
        CSReg_24 <= _GEN_1244;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_25 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h19 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_25 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_25 <= _GEN_281;
      end else begin
        CSReg_25 <= _GEN_1245;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_26 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1a == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_26 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_26 <= _GEN_282;
      end else begin
        CSReg_26 <= _GEN_1246;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_27 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1b == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_27 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_27 <= _GEN_283;
      end else begin
        CSReg_27 <= _GEN_1247;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_28 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1c == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_28 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_28 <= _GEN_284;
      end else begin
        CSReg_28 <= _GEN_1248;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_29 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1d == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_29 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_29 <= _GEN_285;
      end else begin
        CSReg_29 <= _GEN_1249;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_30 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1e == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_30 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_30 <= _GEN_286;
      end else begin
        CSReg_30 <= _GEN_1250;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_31 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h1f == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_31 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_31 <= _GEN_287;
      end else begin
        CSReg_31 <= _GEN_1251;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_32 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h20 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_32 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_32 <= _GEN_288;
      end else begin
        CSReg_32 <= _GEN_1252;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_33 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h21 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_33 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_33 <= _GEN_289;
      end else begin
        CSReg_33 <= _GEN_1253;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_34 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h22 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_34 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_34 <= _GEN_290;
      end else begin
        CSReg_34 <= _GEN_1254;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_35 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h23 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_35 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_35 <= _GEN_291;
      end else begin
        CSReg_35 <= _GEN_1255;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_36 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h24 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_36 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_36 <= _GEN_292;
      end else begin
        CSReg_36 <= _GEN_1256;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_37 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h25 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_37 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_37 <= _GEN_293;
      end else begin
        CSReg_37 <= _GEN_1257;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_38 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h26 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_38 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_38 <= _GEN_294;
      end else begin
        CSReg_38 <= _GEN_1258;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_39 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h27 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_39 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_39 <= _GEN_295;
      end else begin
        CSReg_39 <= _GEN_1259;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_40 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h28 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_40 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_40 <= _GEN_296;
      end else begin
        CSReg_40 <= _GEN_1260;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_41 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h29 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_41 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_41 <= _GEN_297;
      end else begin
        CSReg_41 <= _GEN_1261;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_42 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2a == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_42 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_42 <= _GEN_298;
      end else begin
        CSReg_42 <= _GEN_1262;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_43 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2b == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_43 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_43 <= _GEN_299;
      end else begin
        CSReg_43 <= _GEN_1263;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_44 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2c == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_44 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_44 <= _GEN_300;
      end else begin
        CSReg_44 <= _GEN_1264;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_45 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2d == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_45 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_45 <= _GEN_301;
      end else begin
        CSReg_45 <= _GEN_1265;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_46 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2e == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_46 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_46 <= _GEN_302;
      end else begin
        CSReg_46 <= _GEN_1266;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_47 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h2f == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_47 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_47 <= _GEN_303;
      end else begin
        CSReg_47 <= _GEN_1267;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_48 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h30 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_48 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_48 <= _GEN_304;
      end else begin
        CSReg_48 <= _GEN_1268;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_49 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h31 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_49 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_49 <= _GEN_305;
      end else begin
        CSReg_49 <= _GEN_1269;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_50 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h32 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_50 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_50 <= _GEN_306;
      end else begin
        CSReg_50 <= _GEN_1270;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_51 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h33 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_51 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_51 <= _GEN_307;
      end else begin
        CSReg_51 <= _GEN_1271;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_52 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h34 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_52 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_52 <= _GEN_308;
      end else begin
        CSReg_52 <= _GEN_1272;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_53 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h35 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_53 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_53 <= _GEN_309;
      end else begin
        CSReg_53 <= _GEN_1273;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_54 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h36 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_54 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_54 <= _GEN_310;
      end else begin
        CSReg_54 <= _GEN_1274;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_55 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h37 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_55 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_55 <= _GEN_311;
      end else begin
        CSReg_55 <= _GEN_1275;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_56 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h38 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_56 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_56 <= _GEN_312;
      end else begin
        CSReg_56 <= _GEN_1276;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_57 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h39 == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_57 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_57 <= _GEN_313;
      end else begin
        CSReg_57 <= _GEN_1277;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_58 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3a == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_58 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_58 <= _GEN_314;
      end else begin
        CSReg_58 <= _GEN_1278;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_59 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3b == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_59 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_59 <= _GEN_315;
      end else begin
        CSReg_59 <= _GEN_1279;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_60 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3c == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_60 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_60 <= _GEN_316;
      end else begin
        CSReg_60 <= _GEN_1280;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_61 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3d == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_61 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_61 <= _GEN_317;
      end else begin
        CSReg_61 <= _GEN_1281;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_62 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3e == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_62 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_62 <= _GEN_318;
      end else begin
        CSReg_62 <= _GEN_1282;
      end
    end
    if (reset) begin // @[CSR.scala 23:22]
      CSReg_63 <= 32'h0; // @[CSR.scala 23:22]
    end else if (!(3'h0 == io_CSRType)) begin // @[CSR.scala 27:21]
      if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
        if (6'h3f == io_CSRAddr[5:0]) begin // @[CSR.scala 33:25]
          CSReg_63 <= io_RegFileData; // @[CSR.scala 33:25]
        end
      end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
        CSReg_63 <= _GEN_319;
      end else begin
        CSReg_63 <= _GEN_1283;
      end
    end
    if (reset) begin // @[CSR.scala 25:20]
      out <= 32'h0; // @[CSR.scala 25:20]
    end else if (3'h0 == io_CSRType) begin // @[CSR.scala 27:21]
      out <= 32'h0; // @[CSR.scala 29:11]
    end else if (3'h1 == io_CSRType) begin // @[CSR.scala 27:21]
      out <= _GEN_63; // @[CSR.scala 32:11]
    end else if (3'h2 == io_CSRType) begin // @[CSR.scala 27:21]
      out <= _GEN_63; // @[CSR.scala 36:11]
    end else begin
      out <= _GEN_1219;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  CSReg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  CSReg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  CSReg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  CSReg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  CSReg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  CSReg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  CSReg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  CSReg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  CSReg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  CSReg_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  CSReg_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  CSReg_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  CSReg_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  CSReg_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  CSReg_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  CSReg_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  CSReg_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  CSReg_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  CSReg_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  CSReg_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  CSReg_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  CSReg_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  CSReg_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  CSReg_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  CSReg_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  CSReg_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  CSReg_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  CSReg_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  CSReg_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  CSReg_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  CSReg_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  CSReg_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  CSReg_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  CSReg_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  CSReg_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  CSReg_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  CSReg_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  CSReg_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  CSReg_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  CSReg_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  CSReg_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  CSReg_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  CSReg_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  CSReg_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  CSReg_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  CSReg_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  CSReg_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  CSReg_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  CSReg_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  CSReg_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  CSReg_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  CSReg_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  CSReg_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  CSReg_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  CSReg_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  CSReg_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  CSReg_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  CSReg_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  CSReg_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  CSReg_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  CSReg_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  CSReg_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  CSReg_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  CSReg_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  out = _RAND_64[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rpu_core(
  input         clock,
  input         reset,
  input         io_std_clk,
  input  [31:0] io_boot_addr_0,
  input  [31:0] io_boot_addr_1,
  output [31:0] io_instr_addr,
  input  [31:0] io_instr_data,
  output        io_data_we,
  output [3:0]  io_data_be,
  output [31:0] io_data_addr,
  output [31:0] io_data_wdata,
  input  [31:0] io_data_rdata,
  input         io_IMiss,
  input         io_DMiss
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
`endif // RANDOMIZE_REG_INIT
  wire  tc_clock; // @[rpu_core.scala 103:18]
  wire  tc_reset; // @[rpu_core.scala 103:18]
  wire  tc_io_data_stall; // @[rpu_core.scala 103:18]
  wire  tc_io_control_stall; // @[rpu_core.scala 103:18]
  wire  tc_io_tkend; // @[rpu_core.scala 103:18]
  wire  tc_io_addtk; // @[rpu_core.scala 103:18]
  wire [31:0] tc_io_time; // @[rpu_core.scala 103:18]
  wire [31:0] tc_io_tid; // @[rpu_core.scala 103:18]
  wire [31:0] tc_io_ti; // @[rpu_core.scala 103:18]
  wire  tc_io_wb_pc; // @[rpu_core.scala 103:18]
  wire  tc_io_pc_we; // @[rpu_core.scala 103:18]
  wire  tc_io_ifid_clear; // @[rpu_core.scala 103:18]
  wire  tc_io_ifid_we; // @[rpu_core.scala 103:18]
  wire  tc_io_idex_clear; // @[rpu_core.scala 103:18]
  wire  tc_io_idex_we; // @[rpu_core.scala 103:18]
  wire  tc_io_exmm_clear; // @[rpu_core.scala 103:18]
  wire  tc_io_exmm_we; // @[rpu_core.scala 103:18]
  wire  tc_io_mmwb_clear; // @[rpu_core.scala 103:18]
  wire  tc_io_mmwb_we; // @[rpu_core.scala 103:18]
  wire  tc_io_thread_id_we; // @[rpu_core.scala 103:18]
  wire  tc_io_thread_id_wdata; // @[rpu_core.scala 103:18]
  wire  pcg_clock; // @[rpu_core.scala 105:19]
  wire  pcg_reset; // @[rpu_core.scala 105:19]
  wire [31:0] pcg_io_boot_addr_0; // @[rpu_core.scala 105:19]
  wire [31:0] pcg_io_boot_addr_1; // @[rpu_core.scala 105:19]
  wire  pcg_io_thread_id_we; // @[rpu_core.scala 105:19]
  wire  pcg_io_thread_id_wdata; // @[rpu_core.scala 105:19]
  wire  pcg_io_npc_we; // @[rpu_core.scala 105:19]
  wire [31:0] pcg_io_npc_wdata; // @[rpu_core.scala 105:19]
  wire [31:0] pcg_io_pc; // @[rpu_core.scala 105:19]
  wire  regg_clock; // @[rpu_core.scala 107:20]
  wire  regg_reset; // @[rpu_core.scala 107:20]
  wire  regg_io_TID_Change_En; // @[rpu_core.scala 107:20]
  wire  regg_io_TID_Changed_ID; // @[rpu_core.scala 107:20]
  wire [4:0] regg_io_Raddr1; // @[rpu_core.scala 107:20]
  wire [4:0] regg_io_Raddr2; // @[rpu_core.scala 107:20]
  wire [4:0] regg_io_Raddr3; // @[rpu_core.scala 107:20]
  wire [31:0] regg_io_Rdata1; // @[rpu_core.scala 107:20]
  wire [31:0] regg_io_Rdata2; // @[rpu_core.scala 107:20]
  wire [31:0] regg_io_Rdata3; // @[rpu_core.scala 107:20]
  wire  regg_io_Write_En; // @[rpu_core.scala 107:20]
  wire [4:0] regg_io_Waddr; // @[rpu_core.scala 107:20]
  wire [31:0] regg_io_Wdata; // @[rpu_core.scala 107:20]
  wire [31:0] decoder_io_ir; // @[rpu_core.scala 109:23]
  wire [5:0] decoder_io_instr_type; // @[rpu_core.scala 109:23]
  wire [4:0] decoder_io_rs1; // @[rpu_core.scala 109:23]
  wire [4:0] decoder_io_rs2; // @[rpu_core.scala 109:23]
  wire [4:0] decoder_io_rs3; // @[rpu_core.scala 109:23]
  wire [4:0] decoder_io_rd; // @[rpu_core.scala 109:23]
  wire [31:0] decoder_io_imm; // @[rpu_core.scala 109:23]
  wire [11:0] decoder_io_CSRAddr; // @[rpu_core.scala 109:23]
  wire [5:0] control_io_instr_type; // @[rpu_core.scala 111:23]
  wire  control_io_jump; // @[rpu_core.scala 111:23]
  wire  control_io_branch; // @[rpu_core.scala 111:23]
  wire  control_io_alu_op1_src; // @[rpu_core.scala 111:23]
  wire  control_io_alu_op2_src; // @[rpu_core.scala 111:23]
  wire [3:0] control_io_alu_op; // @[rpu_core.scala 111:23]
  wire [1:0] control_io_alu_result_src; // @[rpu_core.scala 111:23]
  wire [2:0] control_io_comp_op; // @[rpu_core.scala 111:23]
  wire  control_io_r2_src; // @[rpu_core.scala 111:23]
  wire  control_io_tg_we; // @[rpu_core.scala 111:23]
  wire  control_io_ti_we; // @[rpu_core.scala 111:23]
  wire  control_io_to; // @[rpu_core.scala 111:23]
  wire  control_io_addtk; // @[rpu_core.scala 111:23]
  wire  control_io_tkend; // @[rpu_core.scala 111:23]
  wire  control_io_mem_write; // @[rpu_core.scala 111:23]
  wire [3:0] control_io_mem_op; // @[rpu_core.scala 111:23]
  wire  control_io_reg_write; // @[rpu_core.scala 111:23]
  wire [1:0] control_io_reg_write_src; // @[rpu_core.scala 111:23]
  wire [2:0] control_io_csrType; // @[rpu_core.scala 111:23]
  wire [31:0] alu_io_op_a; // @[rpu_core.scala 113:19]
  wire [31:0] alu_io_op_b; // @[rpu_core.scala 113:19]
  wire [31:0] alu_io_csrResult; // @[rpu_core.scala 113:19]
  wire [3:0] alu_io_operation; // @[rpu_core.scala 113:19]
  wire [31:0] alu_io_result; // @[rpu_core.scala 113:19]
  wire [2:0] comp_io_comp_op; // @[rpu_core.scala 115:20]
  wire [31:0] comp_io_op_a; // @[rpu_core.scala 115:20]
  wire [31:0] comp_io_op_b; // @[rpu_core.scala 115:20]
  wire  comp_io_result; // @[rpu_core.scala 115:20]
  wire  tu_clock; // @[rpu_core.scala 117:18]
  wire  tu_reset; // @[rpu_core.scala 117:18]
  wire  tu_io_std_clk; // @[rpu_core.scala 117:18]
  wire  tu_io_ti_we; // @[rpu_core.scala 117:18]
  wire [31:0] tu_io_ti_wdata; // @[rpu_core.scala 117:18]
  wire  tu_io_tg_we; // @[rpu_core.scala 117:18]
  wire [31:0] tu_io_tg_wdata; // @[rpu_core.scala 117:18]
  wire [31:0] tu_io_ti; // @[rpu_core.scala 117:18]
  wire  csr_clock; // @[rpu_core.scala 120:19]
  wire  csr_reset; // @[rpu_core.scala 120:19]
  wire [2:0] csr_io_CSRType; // @[rpu_core.scala 120:19]
  wire [11:0] csr_io_CSRAddr; // @[rpu_core.scala 120:19]
  wire [31:0] csr_io_RegFileData; // @[rpu_core.scala 120:19]
  wire [31:0] csr_io_rsData; // @[rpu_core.scala 120:19]
  wire [31:0] csr_io_CSROut; // @[rpu_core.scala 120:19]
  reg  ifid_stage_regs_valid; // @[rpu_core.scala 129:32]
  reg [31:0] ifid_stage_regs_pc; // @[rpu_core.scala 129:32]
  reg [31:0] ifid_stage_regs_npc; // @[rpu_core.scala 129:32]
  reg [31:0] ifid_stage_regs_ir; // @[rpu_core.scala 129:32]
  reg  idex_stage_regs_valid; // @[rpu_core.scala 164:32]
  reg [31:0] idex_stage_regs_pc; // @[rpu_core.scala 164:32]
  reg [31:0] idex_stage_regs_npc; // @[rpu_core.scala 164:32]
  reg [31:0] idex_stage_regs_r1; // @[rpu_core.scala 164:32]
  reg [31:0] idex_stage_regs_r2; // @[rpu_core.scala 164:32]
  reg [31:0] idex_stage_regs_r3; // @[rpu_core.scala 164:32]
  reg [31:0] idex_stage_regs_imm; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_reg_write; // @[rpu_core.scala 164:32]
  reg [1:0] idex_stage_regs_reg_write_src; // @[rpu_core.scala 164:32]
  reg [4:0] idex_stage_regs_reg_write_addr; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_mem_write; // @[rpu_core.scala 164:32]
  reg [3:0] idex_stage_regs_mem_op; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_jump; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_branch; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_alu_op1_src; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_alu_op2_src; // @[rpu_core.scala 164:32]
  reg [3:0] idex_stage_regs_alu_op; // @[rpu_core.scala 164:32]
  reg [2:0] idex_stage_regs_comp_op; // @[rpu_core.scala 164:32]
  reg [1:0] idex_stage_regs_alu_result_src; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_r2_src; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_tg_we; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_ti_we; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_to; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_addtk; // @[rpu_core.scala 164:32]
  reg  idex_stage_regs_tkend; // @[rpu_core.scala 164:32]
  reg [11:0] idex_stage_regs_csrAddr; // @[rpu_core.scala 164:32]
  reg [2:0] idex_stage_regs_csrType; // @[rpu_core.scala 164:32]
  reg [31:0] exmm_stage_regs_npc; // @[rpu_core.scala 177:32]
  reg [31:0] exmm_stage_regs_alu_result; // @[rpu_core.scala 177:32]
  reg [31:0] exmm_stage_regs_r2; // @[rpu_core.scala 177:32]
  reg  exmm_stage_regs_mem_write; // @[rpu_core.scala 177:32]
  reg [3:0] exmm_stage_regs_mem_op; // @[rpu_core.scala 177:32]
  reg  exmm_stage_regs_reg_write; // @[rpu_core.scala 177:32]
  reg [1:0] exmm_stage_regs_reg_write_src; // @[rpu_core.scala 177:32]
  reg [4:0] exmm_stage_regs_reg_write_addr; // @[rpu_core.scala 177:32]
  reg [31:0] mmwb_stage_regs_npc; // @[rpu_core.scala 188:32]
  reg [31:0] mmwb_stage_regs_alu_result; // @[rpu_core.scala 188:32]
  reg [31:0] mmwb_stage_regs_mem_result; // @[rpu_core.scala 188:32]
  reg  mmwb_stage_regs_reg_write; // @[rpu_core.scala 188:32]
  reg [1:0] mmwb_stage_regs_reg_write_src; // @[rpu_core.scala 188:32]
  reg [4:0] mmwb_stage_regs_reg_write_addr; // @[rpu_core.scala 188:32]
  wire [31:0] _GEN_0 = ifid_stage_regs_valid ? ifid_stage_regs_pc : pcg_io_pc; // @[rpu_core.scala 205:41 206:24 208:24]
  wire [31:0] _GEN_1 = idex_stage_regs_valid ? idex_stage_regs_pc : _GEN_0; // @[rpu_core.scala 203:34 204:24]
  wire  _T = idex_stage_regs_branch & comp_io_result; // @[rpu_core.scala 212:59]
  wire [31:0] _pcg_io_npc_wdata_T_1 = pcg_io_pc + 32'h4; // @[rpu_core.scala 215:37]
  wire [31:0] _GEN_2 = idex_stage_regs_jump | idex_stage_regs_branch & comp_io_result ? alu_io_result :
    _pcg_io_npc_wdata_T_1; // @[rpu_core.scala 212:79 213:24 215:24]
  wire  _GEN_3 = tc_io_pc_we; // @[rpu_core.scala 210:29 211:19 218:19]
  wire [31:0] _GEN_4 = tc_io_pc_we ? _GEN_2 : 32'h0; // @[rpu_core.scala 210:29 219:22]
  wire  _T_4 = ~io_IMiss & ~io_DMiss; // @[rpu_core.scala 227:55]
  wire  _GEN_7 = tc_io_ifid_we & (~io_IMiss & ~io_DMiss) | ifid_stage_regs_valid; // @[rpu_core.scala 227:81 228:27 233:21]
  wire [1:0] _GEN_38 = tc_io_idex_we & _T_4 ? control_io_alu_result_src : 2'h0; // @[rpu_core.scala 154:35 245:81 271:37]
  wire [1:0] idex_stage_reset_alu_result_src = tc_io_idex_clear ? 2'h0 : _GEN_38; // @[rpu_core.scala 243:27 154:35]
  reg [31:0] ts; // @[rpu_core.scala 312:19]
  wire  _data_stall_T_2 = decoder_io_rs1 == idex_stage_regs_reg_write_addr; // @[rpu_core.scala 323:35]
  wire  _data_stall_T_3 = idex_stage_regs_reg_write & idex_stage_regs_reg_write_addr != 5'h0 & _data_stall_T_2; // @[rpu_core.scala 322:86]
  wire  _data_stall_T_4 = decoder_io_rs2 == idex_stage_regs_reg_write_addr; // @[rpu_core.scala 324:35]
  wire  _data_stall_T_5 = _data_stall_T_3 | _data_stall_T_4; // @[rpu_core.scala 323:71]
  wire  _data_stall_T_6 = decoder_io_rs3 == idex_stage_regs_reg_write_addr; // @[rpu_core.scala 325:35]
  wire  _data_stall_T_7 = _data_stall_T_5 | _data_stall_T_6; // @[rpu_core.scala 324:71]
  wire  _data_stall_T_10 = decoder_io_rs1 == exmm_stage_regs_reg_write_addr; // @[rpu_core.scala 327:35]
  wire  _data_stall_T_11 = exmm_stage_regs_reg_write & exmm_stage_regs_reg_write_addr != 5'h0 & _data_stall_T_10; // @[rpu_core.scala 326:86]
  wire  _data_stall_T_12 = decoder_io_rs2 == exmm_stage_regs_reg_write_addr; // @[rpu_core.scala 328:35]
  wire  _data_stall_T_13 = _data_stall_T_11 | _data_stall_T_12; // @[rpu_core.scala 327:71]
  wire  _data_stall_T_14 = decoder_io_rs3 == exmm_stage_regs_reg_write_addr; // @[rpu_core.scala 329:35]
  wire  _data_stall_T_15 = _data_stall_T_13 | _data_stall_T_14; // @[rpu_core.scala 328:71]
  wire  _data_stall_T_16 = _data_stall_T_7 | _data_stall_T_15; // @[rpu_core.scala 325:72]
  wire  _data_stall_T_19 = decoder_io_rs1 == mmwb_stage_regs_reg_write_addr; // @[rpu_core.scala 331:35]
  wire  _data_stall_T_20 = mmwb_stage_regs_reg_write & mmwb_stage_regs_reg_write_addr != 5'h0 & _data_stall_T_19; // @[rpu_core.scala 330:86]
  wire  _data_stall_T_21 = decoder_io_rs2 == mmwb_stage_regs_reg_write_addr; // @[rpu_core.scala 332:35]
  wire  _data_stall_T_22 = _data_stall_T_20 | _data_stall_T_21; // @[rpu_core.scala 331:71]
  wire  _data_stall_T_23 = decoder_io_rs3 == mmwb_stage_regs_reg_write_addr; // @[rpu_core.scala 333:35]
  wire  _data_stall_T_24 = _data_stall_T_22 | _data_stall_T_23; // @[rpu_core.scala 332:71]
  wire [31:0] _GEN_80 = 2'h2 == idex_stage_regs_alu_result_src ? tu_io_ti : exmm_stage_regs_alu_result; // @[rpu_core.scala 177:32 354:45 362:36]
  wire [31:0] _GEN_81 = 2'h1 == idex_stage_regs_alu_result_src ? ts : _GEN_80; // @[rpu_core.scala 354:45 359:36]
  wire [31:0] _io_data_addr_T_1 = {exmm_stage_regs_alu_result[31:2],2'h0}; // @[Cat.scala 31:58]
  wire [6:0] _io_data_be_T_1 = 7'h1 << exmm_stage_regs_alu_result[1:0]; // @[rpu_core.scala 390:32]
  wire [3:0] _GEN_102 = exmm_stage_regs_alu_result[1] ? 4'hc : 4'h3; // @[rpu_core.scala 394:46 395:22 397:22]
  wire [31:0] _GEN_103 = 4'h8 == exmm_stage_regs_mem_op ? _io_data_addr_T_1 : 32'h0; // @[rpu_core.scala 385:18 387:37 401:22]
  wire [3:0] _GEN_104 = 4'h8 == exmm_stage_regs_mem_op ? 4'hf : 4'h0; // @[rpu_core.scala 386:16 387:37 402:20]
  wire [31:0] _GEN_105 = 4'h7 == exmm_stage_regs_mem_op ? _io_data_addr_T_1 : _GEN_103; // @[rpu_core.scala 387:37 393:22]
  wire [3:0] _GEN_106 = 4'h7 == exmm_stage_regs_mem_op ? _GEN_102 : _GEN_104; // @[rpu_core.scala 387:37]
  wire [31:0] _GEN_107 = 4'h6 == exmm_stage_regs_mem_op ? _io_data_addr_T_1 : _GEN_105; // @[rpu_core.scala 387:37 389:22]
  wire [6:0] _GEN_108 = 4'h6 == exmm_stage_regs_mem_op ? _io_data_be_T_1 : {{3'd0}, _GEN_106}; // @[rpu_core.scala 387:37 390:20]
  wire [6:0] _GEN_112 = exmm_stage_regs_mem_write ? _GEN_108 : 7'h0; // @[rpu_core.scala 382:36 408:16]
  wire [23:0] _mmwb_stage_regs_mem_result_T_2 = io_data_rdata[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _mmwb_stage_regs_mem_result_T_4 = {_mmwb_stage_regs_mem_result_T_2,io_data_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _mmwb_stage_regs_mem_result_T_6 = {24'h0,io_data_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [15:0] _mmwb_stage_regs_mem_result_T_9 = io_data_rdata[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _mmwb_stage_regs_mem_result_T_11 = {_mmwb_stage_regs_mem_result_T_9,io_data_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _mmwb_stage_regs_mem_result_T_13 = {16'h0,io_data_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_113 = 4'h3 == exmm_stage_regs_mem_op ? io_data_rdata : 32'h0; // @[rpu_core.scala 418:32 419:37 433:36]
  wire [31:0] _GEN_114 = 4'h5 == exmm_stage_regs_mem_op ? _mmwb_stage_regs_mem_result_T_13 : _GEN_113; // @[rpu_core.scala 419:37 430:36]
  wire [31:0] _GEN_115 = 4'h2 == exmm_stage_regs_mem_op ? _mmwb_stage_regs_mem_result_T_11 : _GEN_114; // @[rpu_core.scala 419:37 427:36]
  wire [31:0] _GEN_116 = 4'h4 == exmm_stage_regs_mem_op ? _mmwb_stage_regs_mem_result_T_6 : _GEN_115; // @[rpu_core.scala 419:37 424:36]
  wire [31:0] _GEN_133 = 2'h1 == mmwb_stage_regs_reg_write_src ? mmwb_stage_regs_alu_result : mmwb_stage_regs_npc; // @[rpu_core.scala 447:43 452:23]
  wire [31:0] _GEN_134 = 2'h0 == mmwb_stage_regs_reg_write_src ? mmwb_stage_regs_mem_result : _GEN_133; // @[rpu_core.scala 447:43 449:23]
  rpu_thread_control tc ( // @[rpu_core.scala 103:18]
    .clock(tc_clock),
    .reset(tc_reset),
    .io_data_stall(tc_io_data_stall),
    .io_control_stall(tc_io_control_stall),
    .io_tkend(tc_io_tkend),
    .io_addtk(tc_io_addtk),
    .io_time(tc_io_time),
    .io_tid(tc_io_tid),
    .io_ti(tc_io_ti),
    .io_wb_pc(tc_io_wb_pc),
    .io_pc_we(tc_io_pc_we),
    .io_ifid_clear(tc_io_ifid_clear),
    .io_ifid_we(tc_io_ifid_we),
    .io_idex_clear(tc_io_idex_clear),
    .io_idex_we(tc_io_idex_we),
    .io_exmm_clear(tc_io_exmm_clear),
    .io_exmm_we(tc_io_exmm_we),
    .io_mmwb_clear(tc_io_mmwb_clear),
    .io_mmwb_we(tc_io_mmwb_we),
    .io_thread_id_we(tc_io_thread_id_we),
    .io_thread_id_wdata(tc_io_thread_id_wdata)
  );
  rpu_pc_group pcg ( // @[rpu_core.scala 105:19]
    .clock(pcg_clock),
    .reset(pcg_reset),
    .io_boot_addr_0(pcg_io_boot_addr_0),
    .io_boot_addr_1(pcg_io_boot_addr_1),
    .io_thread_id_we(pcg_io_thread_id_we),
    .io_thread_id_wdata(pcg_io_thread_id_wdata),
    .io_npc_we(pcg_io_npc_we),
    .io_npc_wdata(pcg_io_npc_wdata),
    .io_pc(pcg_io_pc)
  );
  RegisterFileGroup regg ( // @[rpu_core.scala 107:20]
    .clock(regg_clock),
    .reset(regg_reset),
    .io_TID_Change_En(regg_io_TID_Change_En),
    .io_TID_Changed_ID(regg_io_TID_Changed_ID),
    .io_Raddr1(regg_io_Raddr1),
    .io_Raddr2(regg_io_Raddr2),
    .io_Raddr3(regg_io_Raddr3),
    .io_Rdata1(regg_io_Rdata1),
    .io_Rdata2(regg_io_Rdata2),
    .io_Rdata3(regg_io_Rdata3),
    .io_Write_En(regg_io_Write_En),
    .io_Waddr(regg_io_Waddr),
    .io_Wdata(regg_io_Wdata)
  );
  rpu_decoder decoder ( // @[rpu_core.scala 109:23]
    .io_ir(decoder_io_ir),
    .io_instr_type(decoder_io_instr_type),
    .io_rs1(decoder_io_rs1),
    .io_rs2(decoder_io_rs2),
    .io_rs3(decoder_io_rs3),
    .io_rd(decoder_io_rd),
    .io_imm(decoder_io_imm),
    .io_CSRAddr(decoder_io_CSRAddr)
  );
  rpu_control control ( // @[rpu_core.scala 111:23]
    .io_instr_type(control_io_instr_type),
    .io_jump(control_io_jump),
    .io_branch(control_io_branch),
    .io_alu_op1_src(control_io_alu_op1_src),
    .io_alu_op2_src(control_io_alu_op2_src),
    .io_alu_op(control_io_alu_op),
    .io_alu_result_src(control_io_alu_result_src),
    .io_comp_op(control_io_comp_op),
    .io_r2_src(control_io_r2_src),
    .io_tg_we(control_io_tg_we),
    .io_ti_we(control_io_ti_we),
    .io_to(control_io_to),
    .io_addtk(control_io_addtk),
    .io_tkend(control_io_tkend),
    .io_mem_write(control_io_mem_write),
    .io_mem_op(control_io_mem_op),
    .io_reg_write(control_io_reg_write),
    .io_reg_write_src(control_io_reg_write_src),
    .io_csrType(control_io_csrType)
  );
  rpu_alu alu ( // @[rpu_core.scala 113:19]
    .io_op_a(alu_io_op_a),
    .io_op_b(alu_io_op_b),
    .io_csrResult(alu_io_csrResult),
    .io_operation(alu_io_operation),
    .io_result(alu_io_result)
  );
  rpu_comp comp ( // @[rpu_core.scala 115:20]
    .io_comp_op(comp_io_comp_op),
    .io_op_a(comp_io_op_a),
    .io_op_b(comp_io_op_b),
    .io_result(comp_io_result)
  );
  rpu_time_unit tu ( // @[rpu_core.scala 117:18]
    .clock(tu_clock),
    .reset(tu_reset),
    .io_std_clk(tu_io_std_clk),
    .io_ti_we(tu_io_ti_we),
    .io_ti_wdata(tu_io_ti_wdata),
    .io_tg_we(tu_io_tg_we),
    .io_tg_wdata(tu_io_tg_wdata),
    .io_ti(tu_io_ti)
  );
  CSR csr ( // @[rpu_core.scala 120:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_CSRType(csr_io_CSRType),
    .io_CSRAddr(csr_io_CSRAddr),
    .io_RegFileData(csr_io_RegFileData),
    .io_rsData(csr_io_rsData),
    .io_CSROut(csr_io_CSROut)
  );
  assign io_instr_addr = pcg_io_pc; // @[rpu_core.scala 223:17]
  assign io_data_we = exmm_stage_regs_mem_write; // @[rpu_core.scala 382:36 383:16 406:16]
  assign io_data_be = _GEN_112[3:0];
  assign io_data_addr = exmm_stage_regs_mem_write ? _GEN_107 : _io_data_addr_T_1; // @[rpu_core.scala 382:36 409:18]
  assign io_data_wdata = exmm_stage_regs_mem_write ? exmm_stage_regs_r2 : 32'h0; // @[rpu_core.scala 382:36 384:19 407:19]
  assign tc_clock = clock;
  assign tc_reset = reset;
  assign tc_io_data_stall = _data_stall_T_16 | _data_stall_T_24; // @[rpu_core.scala 329:72]
  assign tc_io_control_stall = idex_stage_regs_jump | _T; // @[rpu_core.scala 335:41]
  assign tc_io_tkend = idex_stage_regs_tkend; // @[rpu_core.scala 342:15]
  assign tc_io_addtk = idex_stage_regs_addtk; // @[rpu_core.scala 343:15]
  assign tc_io_time = idex_stage_regs_r1; // @[rpu_core.scala 344:14]
  assign tc_io_tid = idex_stage_regs_r2; // @[rpu_core.scala 345:13]
  assign tc_io_ti = tu_io_ti; // @[rpu_core.scala 337:12]
  assign pcg_clock = clock;
  assign pcg_reset = reset;
  assign pcg_io_boot_addr_0 = io_boot_addr_0; // @[rpu_core.scala 192:20]
  assign pcg_io_boot_addr_1 = io_boot_addr_1; // @[rpu_core.scala 192:20]
  assign pcg_io_thread_id_we = tc_io_thread_id_we; // @[rpu_core.scala 195:23]
  assign pcg_io_thread_id_wdata = tc_io_thread_id_wdata; // @[rpu_core.scala 196:26]
  assign pcg_io_npc_we = tc_io_wb_pc | _GEN_3; // @[rpu_core.scala 201:22 202:19]
  assign pcg_io_npc_wdata = tc_io_wb_pc ? _GEN_1 : _GEN_4; // @[rpu_core.scala 201:22]
  assign regg_clock = clock;
  assign regg_reset = reset;
  assign regg_io_TID_Change_En = tc_io_thread_id_we; // @[rpu_core.scala 197:25]
  assign regg_io_TID_Changed_ID = tc_io_thread_id_wdata; // @[rpu_core.scala 198:26]
  assign regg_io_Raddr1 = decoder_io_rs1; // @[rpu_core.scala 239:18]
  assign regg_io_Raddr2 = decoder_io_rs2; // @[rpu_core.scala 240:18]
  assign regg_io_Raddr3 = decoder_io_rs3; // @[rpu_core.scala 241:18]
  assign regg_io_Write_En = mmwb_stage_regs_reg_write; // @[rpu_core.scala 443:20]
  assign regg_io_Waddr = mmwb_stage_regs_reg_write_addr; // @[rpu_core.scala 444:17]
  assign regg_io_Wdata = mmwb_stage_regs_reg_write ? _GEN_134 : mmwb_stage_regs_npc; // @[rpu_core.scala 445:17 446:36]
  assign decoder_io_ir = ifid_stage_regs_ir; // @[rpu_core.scala 237:17]
  assign control_io_instr_type = decoder_io_instr_type; // @[rpu_core.scala 238:25]
  assign alu_io_op_a = idex_stage_regs_alu_op1_src ? idex_stage_regs_pc : idex_stage_regs_r1; // @[rpu_core.scala 292:59 293:17 295:17]
  assign alu_io_op_b = idex_stage_regs_alu_op2_src ? idex_stage_regs_imm : idex_stage_regs_r2; // @[rpu_core.scala 297:60 298:17 300:17]
  assign alu_io_csrResult = csr_io_CSROut; // @[rpu_core.scala 304:20]
  assign alu_io_operation = idex_stage_regs_alu_op; // @[rpu_core.scala 302:20]
  assign comp_io_comp_op = idex_stage_regs_comp_op; // @[rpu_core.scala 290:19]
  assign comp_io_op_a = idex_stage_regs_r1; // @[rpu_core.scala 288:16]
  assign comp_io_op_b = idex_stage_regs_r2; // @[rpu_core.scala 289:16]
  assign tu_clock = clock;
  assign tu_reset = reset;
  assign tu_io_std_clk = io_std_clk; // @[rpu_core.scala 306:17]
  assign tu_io_ti_we = idex_stage_regs_ti_we; // @[rpu_core.scala 307:15]
  assign tu_io_ti_wdata = idex_stage_regs_r1; // @[rpu_core.scala 308:18]
  assign tu_io_tg_we = idex_stage_regs_tg_we; // @[rpu_core.scala 309:15]
  assign tu_io_tg_wdata = idex_stage_regs_r1; // @[rpu_core.scala 310:18]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_CSRType = idex_stage_regs_csrType; // @[rpu_core.scala 284:18]
  assign csr_io_CSRAddr = idex_stage_regs_csrAddr; // @[rpu_core.scala 283:18]
  assign csr_io_RegFileData = idex_stage_regs_r1; // @[rpu_core.scala 286:22]
  assign csr_io_rsData = idex_stage_regs_imm; // @[rpu_core.scala 285:17]
  always @(posedge clock) begin
    if (reset) begin // @[rpu_core.scala 129:32]
      ifid_stage_regs_valid <= 1'h0; // @[rpu_core.scala 129:32]
    end else if (tc_io_ifid_clear) begin // @[rpu_core.scala 225:27]
      ifid_stage_regs_valid <= 1'h0; // @[rpu_core.scala 226:21]
    end else begin
      ifid_stage_regs_valid <= _GEN_7;
    end
    if (reset) begin // @[rpu_core.scala 129:32]
      ifid_stage_regs_pc <= 32'h0; // @[rpu_core.scala 129:32]
    end else if (tc_io_ifid_clear) begin // @[rpu_core.scala 225:27]
      ifid_stage_regs_pc <= 32'h0; // @[rpu_core.scala 226:21]
    end else if (tc_io_ifid_we & (~io_IMiss & ~io_DMiss)) begin // @[rpu_core.scala 227:81]
      ifid_stage_regs_pc <= pcg_io_pc; // @[rpu_core.scala 229:24]
    end
    if (reset) begin // @[rpu_core.scala 129:32]
      ifid_stage_regs_npc <= 32'h0; // @[rpu_core.scala 129:32]
    end else if (tc_io_ifid_clear) begin // @[rpu_core.scala 225:27]
      ifid_stage_regs_npc <= 32'h0; // @[rpu_core.scala 226:21]
    end else if (tc_io_ifid_we & (~io_IMiss & ~io_DMiss)) begin // @[rpu_core.scala 227:81]
      ifid_stage_regs_npc <= _pcg_io_npc_wdata_T_1; // @[rpu_core.scala 230:25]
    end
    if (reset) begin // @[rpu_core.scala 129:32]
      ifid_stage_regs_ir <= 32'h0; // @[rpu_core.scala 129:32]
    end else if (tc_io_ifid_clear) begin // @[rpu_core.scala 225:27]
      ifid_stage_regs_ir <= 32'h0; // @[rpu_core.scala 226:21]
    end else if (tc_io_ifid_we & (~io_IMiss & ~io_DMiss)) begin // @[rpu_core.scala 227:81]
      ifid_stage_regs_ir <= io_instr_data; // @[rpu_core.scala 231:24]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_valid <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_valid <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_valid <= ifid_stage_regs_valid; // @[rpu_core.scala 246:27]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_pc <= 32'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_pc <= 32'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_pc <= ifid_stage_regs_pc; // @[rpu_core.scala 247:24]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_npc <= 32'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_npc <= 32'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_npc <= ifid_stage_regs_npc; // @[rpu_core.scala 248:25]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_r1 <= 32'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_r1 <= 32'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_r1 <= regg_io_Rdata1; // @[rpu_core.scala 249:24]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_r2 <= 32'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_r2 <= 32'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_r2 <= regg_io_Rdata2; // @[rpu_core.scala 250:24]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_r3 <= 32'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_r3 <= 32'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_r3 <= regg_io_Rdata3; // @[rpu_core.scala 251:24]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_imm <= 32'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_imm <= 32'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_imm <= decoder_io_imm; // @[rpu_core.scala 252:25]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_reg_write <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_reg_write <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_reg_write <= control_io_reg_write; // @[rpu_core.scala 260:31]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_reg_write_src <= 2'h1; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_reg_write_src <= 2'h1; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_reg_write_src <= control_io_reg_write_src; // @[rpu_core.scala 261:35]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_reg_write_addr <= 5'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_reg_write_addr <= 5'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_reg_write_addr <= decoder_io_rd; // @[rpu_core.scala 262:36]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_mem_write <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_mem_write <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_mem_write <= control_io_mem_write; // @[rpu_core.scala 263:31]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_mem_op <= 4'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_mem_op <= 4'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_mem_op <= control_io_mem_op; // @[rpu_core.scala 264:28]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_jump <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_jump <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_jump <= control_io_jump; // @[rpu_core.scala 265:26]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_branch <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_branch <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_branch <= control_io_branch; // @[rpu_core.scala 266:28]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_alu_op1_src <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_alu_op1_src <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_alu_op1_src <= control_io_alu_op1_src; // @[rpu_core.scala 267:33]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_alu_op2_src <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_alu_op2_src <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_alu_op2_src <= control_io_alu_op2_src; // @[rpu_core.scala 268:33]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_alu_op <= 4'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_alu_op <= 4'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_alu_op <= control_io_alu_op; // @[rpu_core.scala 269:28]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_comp_op <= 3'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_comp_op <= 3'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_comp_op <= control_io_comp_op; // @[rpu_core.scala 270:29]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_alu_result_src <= idex_stage_reset_alu_result_src; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_alu_result_src <= idex_stage_reset_alu_result_src; // @[rpu_core.scala 244:21]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_r2_src <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_r2_src <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_r2_src <= control_io_r2_src; // @[rpu_core.scala 272:28]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_tg_we <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_tg_we <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_tg_we <= control_io_tg_we; // @[rpu_core.scala 273:27]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_ti_we <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_ti_we <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_ti_we <= control_io_ti_we; // @[rpu_core.scala 274:27]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_to <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_to <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_to <= control_io_to; // @[rpu_core.scala 275:24]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_addtk <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_addtk <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_addtk <= control_io_addtk; // @[rpu_core.scala 276:27]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_tkend <= 1'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_tkend <= 1'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_tkend <= control_io_tkend; // @[rpu_core.scala 277:27]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_csrAddr <= 12'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_csrAddr <= 12'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_csrAddr <= decoder_io_CSRAddr; // @[rpu_core.scala 258:29]
    end
    if (reset) begin // @[rpu_core.scala 164:32]
      idex_stage_regs_csrType <= 3'h0; // @[rpu_core.scala 164:32]
    end else if (tc_io_idex_clear) begin // @[rpu_core.scala 243:27]
      idex_stage_regs_csrType <= 3'h0; // @[rpu_core.scala 244:21]
    end else if (tc_io_idex_we & _T_4) begin // @[rpu_core.scala 245:81]
      idex_stage_regs_csrType <= control_io_csrType; // @[rpu_core.scala 257:29]
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_npc <= 32'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_npc <= 32'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      exmm_stage_regs_npc <= idex_stage_regs_npc; // @[rpu_core.scala 353:25]
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_alu_result <= 32'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_alu_result <= 32'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      if (2'h0 == idex_stage_regs_alu_result_src) begin // @[rpu_core.scala 354:45]
        exmm_stage_regs_alu_result <= alu_io_result; // @[rpu_core.scala 356:36]
      end else begin
        exmm_stage_regs_alu_result <= _GEN_81;
      end
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_r2 <= 32'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_r2 <= 32'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      if (idex_stage_regs_r2_src) begin // @[rpu_core.scala 365:51]
        exmm_stage_regs_r2 <= idex_stage_regs_r3; // @[rpu_core.scala 366:26]
      end else begin
        exmm_stage_regs_r2 <= idex_stage_regs_r2; // @[rpu_core.scala 368:26]
      end
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_mem_write <= 1'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_mem_write <= 1'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      exmm_stage_regs_mem_write <= idex_stage_regs_mem_write; // @[rpu_core.scala 370:31]
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_mem_op <= 4'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_mem_op <= 4'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      exmm_stage_regs_mem_op <= idex_stage_regs_mem_op; // @[rpu_core.scala 371:28]
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_reg_write <= 1'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_reg_write <= 1'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      exmm_stage_regs_reg_write <= idex_stage_regs_reg_write; // @[rpu_core.scala 372:31]
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_reg_write_src <= 2'h1; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_reg_write_src <= 2'h1; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      exmm_stage_regs_reg_write_src <= idex_stage_regs_reg_write_src; // @[rpu_core.scala 373:35]
    end
    if (reset) begin // @[rpu_core.scala 177:32]
      exmm_stage_regs_reg_write_addr <= 5'h0; // @[rpu_core.scala 177:32]
    end else if (tc_io_exmm_clear) begin // @[rpu_core.scala 349:27]
      exmm_stage_regs_reg_write_addr <= 5'h0; // @[rpu_core.scala 350:21]
    end else if (tc_io_exmm_we & _T_4) begin // @[rpu_core.scala 351:81]
      exmm_stage_regs_reg_write_addr <= idex_stage_regs_reg_write_addr; // @[rpu_core.scala 374:36]
    end
    if (reset) begin // @[rpu_core.scala 188:32]
      mmwb_stage_regs_npc <= 32'h0; // @[rpu_core.scala 188:32]
    end else if (tc_io_mmwb_clear) begin // @[rpu_core.scala 412:27]
      mmwb_stage_regs_npc <= 32'h0; // @[rpu_core.scala 413:21]
    end else if (tc_io_mmwb_we & _T_4) begin // @[rpu_core.scala 414:81]
      mmwb_stage_regs_npc <= exmm_stage_regs_npc; // @[rpu_core.scala 416:25]
    end
    if (reset) begin // @[rpu_core.scala 188:32]
      mmwb_stage_regs_alu_result <= 32'h0; // @[rpu_core.scala 188:32]
    end else if (tc_io_mmwb_clear) begin // @[rpu_core.scala 412:27]
      mmwb_stage_regs_alu_result <= 32'h0; // @[rpu_core.scala 413:21]
    end else if (tc_io_mmwb_we & _T_4) begin // @[rpu_core.scala 414:81]
      mmwb_stage_regs_alu_result <= exmm_stage_regs_alu_result; // @[rpu_core.scala 417:32]
    end
    if (reset) begin // @[rpu_core.scala 188:32]
      mmwb_stage_regs_mem_result <= 32'h0; // @[rpu_core.scala 188:32]
    end else if (tc_io_mmwb_clear) begin // @[rpu_core.scala 412:27]
      mmwb_stage_regs_mem_result <= 32'h0; // @[rpu_core.scala 413:21]
    end else if (tc_io_mmwb_we & _T_4) begin // @[rpu_core.scala 414:81]
      if (4'h1 == exmm_stage_regs_mem_op) begin // @[rpu_core.scala 419:37]
        mmwb_stage_regs_mem_result <= _mmwb_stage_regs_mem_result_T_4; // @[rpu_core.scala 421:36]
      end else begin
        mmwb_stage_regs_mem_result <= _GEN_116;
      end
    end
    if (reset) begin // @[rpu_core.scala 188:32]
      mmwb_stage_regs_reg_write <= 1'h0; // @[rpu_core.scala 188:32]
    end else if (tc_io_mmwb_clear) begin // @[rpu_core.scala 412:27]
      mmwb_stage_regs_reg_write <= 1'h0; // @[rpu_core.scala 413:21]
    end else if (tc_io_mmwb_we & _T_4) begin // @[rpu_core.scala 414:81]
      mmwb_stage_regs_reg_write <= exmm_stage_regs_reg_write; // @[rpu_core.scala 436:31]
    end
    if (reset) begin // @[rpu_core.scala 188:32]
      mmwb_stage_regs_reg_write_src <= 2'h1; // @[rpu_core.scala 188:32]
    end else if (tc_io_mmwb_clear) begin // @[rpu_core.scala 412:27]
      mmwb_stage_regs_reg_write_src <= 2'h1; // @[rpu_core.scala 413:21]
    end else if (tc_io_mmwb_we & _T_4) begin // @[rpu_core.scala 414:81]
      mmwb_stage_regs_reg_write_src <= exmm_stage_regs_reg_write_src; // @[rpu_core.scala 437:35]
    end
    if (reset) begin // @[rpu_core.scala 188:32]
      mmwb_stage_regs_reg_write_addr <= 5'h0; // @[rpu_core.scala 188:32]
    end else if (tc_io_mmwb_clear) begin // @[rpu_core.scala 412:27]
      mmwb_stage_regs_reg_write_addr <= 5'h0; // @[rpu_core.scala 413:21]
    end else if (tc_io_mmwb_we & _T_4) begin // @[rpu_core.scala 414:81]
      mmwb_stage_regs_reg_write_addr <= exmm_stage_regs_reg_write_addr; // @[rpu_core.scala 438:36]
    end
    if (reset) begin // @[rpu_core.scala 312:19]
      ts <= 32'h0; // @[rpu_core.scala 312:19]
    end else if (idex_stage_regs_to & tc_io_exmm_we) begin // @[rpu_core.scala 313:46]
      ts <= tu_io_ti; // @[rpu_core.scala 314:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ifid_stage_regs_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifid_stage_regs_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ifid_stage_regs_npc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ifid_stage_regs_ir = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  idex_stage_regs_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  idex_stage_regs_pc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  idex_stage_regs_npc = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  idex_stage_regs_r1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  idex_stage_regs_r2 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  idex_stage_regs_r3 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  idex_stage_regs_imm = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  idex_stage_regs_reg_write = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  idex_stage_regs_reg_write_src = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  idex_stage_regs_reg_write_addr = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  idex_stage_regs_mem_write = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  idex_stage_regs_mem_op = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  idex_stage_regs_jump = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  idex_stage_regs_branch = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  idex_stage_regs_alu_op1_src = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  idex_stage_regs_alu_op2_src = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  idex_stage_regs_alu_op = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  idex_stage_regs_comp_op = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  idex_stage_regs_alu_result_src = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  idex_stage_regs_r2_src = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  idex_stage_regs_tg_we = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  idex_stage_regs_ti_we = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  idex_stage_regs_to = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  idex_stage_regs_addtk = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  idex_stage_regs_tkend = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  idex_stage_regs_csrAddr = _RAND_29[11:0];
  _RAND_30 = {1{`RANDOM}};
  idex_stage_regs_csrType = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  exmm_stage_regs_npc = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  exmm_stage_regs_alu_result = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  exmm_stage_regs_r2 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  exmm_stage_regs_mem_write = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  exmm_stage_regs_mem_op = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  exmm_stage_regs_reg_write = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  exmm_stage_regs_reg_write_src = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  exmm_stage_regs_reg_write_addr = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  mmwb_stage_regs_npc = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mmwb_stage_regs_alu_result = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mmwb_stage_regs_mem_result = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mmwb_stage_regs_reg_write = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  mmwb_stage_regs_reg_write_src = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  mmwb_stage_regs_reg_write_addr = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  ts = _RAND_45[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache(
  input         clock,
  input         reset,
  input  [31:0] io_addr,
  input         io_r_req,
  input         io_w_req,
  input  [31:0] io_writedata,
  input  [3:0]  io_writeMask,
  output [31:0] io_outdata,
  output        io_miss,
  output [8:0]  io_mem_addr,
  output        io_mem_rd_req,
  output        io_mem_wr_req,
  output [31:0] io_mem_wr_line_0,
  output [31:0] io_mem_wr_line_1,
  output [31:0] io_mem_wr_line_2,
  output [31:0] io_mem_wr_line_3,
  output [31:0] io_mem_wr_line_4,
  output [31:0] io_mem_wr_line_5,
  output [31:0] io_mem_wr_line_6,
  output [31:0] io_mem_wr_line_7,
  input  [31:0] io_mem_rd_line_0,
  input  [31:0] io_mem_rd_line_1,
  input  [31:0] io_mem_rd_line_2,
  input  [31:0] io_mem_rd_line_3,
  input  [31:0] io_mem_rd_line_4,
  input  [31:0] io_mem_rd_line_5,
  input  [31:0] io_mem_rd_line_6,
  input  [31:0] io_mem_rd_line_7,
  input         io_cacheAXI_gnt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] CacheMem_0_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_0_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_1_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_2_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_3_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_4_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_5_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_6_7_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_0_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_1_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_2_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_3_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_4_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_5_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_6_7; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_0; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_1; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_2; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_3; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_4; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_5; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_6; // @[Cache.scala 53:25]
  reg [31:0] CacheMem_7_7_7; // @[Cache.scala 53:25]
  reg [5:0] cache_tags_0_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_0_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_1_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_2_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_3_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_4_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_5_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_6_7; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_0; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_1; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_2; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_3; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_4; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_5; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_6; // @[Cache.scala 56:27]
  reg [5:0] cache_tags_7_7; // @[Cache.scala 56:27]
  reg  valid_0_0; // @[Cache.scala 57:22]
  reg  valid_0_1; // @[Cache.scala 57:22]
  reg  valid_0_2; // @[Cache.scala 57:22]
  reg  valid_0_3; // @[Cache.scala 57:22]
  reg  valid_0_4; // @[Cache.scala 57:22]
  reg  valid_0_5; // @[Cache.scala 57:22]
  reg  valid_0_6; // @[Cache.scala 57:22]
  reg  valid_0_7; // @[Cache.scala 57:22]
  reg  valid_1_0; // @[Cache.scala 57:22]
  reg  valid_1_1; // @[Cache.scala 57:22]
  reg  valid_1_2; // @[Cache.scala 57:22]
  reg  valid_1_3; // @[Cache.scala 57:22]
  reg  valid_1_4; // @[Cache.scala 57:22]
  reg  valid_1_5; // @[Cache.scala 57:22]
  reg  valid_1_6; // @[Cache.scala 57:22]
  reg  valid_1_7; // @[Cache.scala 57:22]
  reg  valid_2_0; // @[Cache.scala 57:22]
  reg  valid_2_1; // @[Cache.scala 57:22]
  reg  valid_2_2; // @[Cache.scala 57:22]
  reg  valid_2_3; // @[Cache.scala 57:22]
  reg  valid_2_4; // @[Cache.scala 57:22]
  reg  valid_2_5; // @[Cache.scala 57:22]
  reg  valid_2_6; // @[Cache.scala 57:22]
  reg  valid_2_7; // @[Cache.scala 57:22]
  reg  valid_3_0; // @[Cache.scala 57:22]
  reg  valid_3_1; // @[Cache.scala 57:22]
  reg  valid_3_2; // @[Cache.scala 57:22]
  reg  valid_3_3; // @[Cache.scala 57:22]
  reg  valid_3_4; // @[Cache.scala 57:22]
  reg  valid_3_5; // @[Cache.scala 57:22]
  reg  valid_3_6; // @[Cache.scala 57:22]
  reg  valid_3_7; // @[Cache.scala 57:22]
  reg  valid_4_0; // @[Cache.scala 57:22]
  reg  valid_4_1; // @[Cache.scala 57:22]
  reg  valid_4_2; // @[Cache.scala 57:22]
  reg  valid_4_3; // @[Cache.scala 57:22]
  reg  valid_4_4; // @[Cache.scala 57:22]
  reg  valid_4_5; // @[Cache.scala 57:22]
  reg  valid_4_6; // @[Cache.scala 57:22]
  reg  valid_4_7; // @[Cache.scala 57:22]
  reg  valid_5_0; // @[Cache.scala 57:22]
  reg  valid_5_1; // @[Cache.scala 57:22]
  reg  valid_5_2; // @[Cache.scala 57:22]
  reg  valid_5_3; // @[Cache.scala 57:22]
  reg  valid_5_4; // @[Cache.scala 57:22]
  reg  valid_5_5; // @[Cache.scala 57:22]
  reg  valid_5_6; // @[Cache.scala 57:22]
  reg  valid_5_7; // @[Cache.scala 57:22]
  reg  valid_6_0; // @[Cache.scala 57:22]
  reg  valid_6_1; // @[Cache.scala 57:22]
  reg  valid_6_2; // @[Cache.scala 57:22]
  reg  valid_6_3; // @[Cache.scala 57:22]
  reg  valid_6_4; // @[Cache.scala 57:22]
  reg  valid_6_5; // @[Cache.scala 57:22]
  reg  valid_6_6; // @[Cache.scala 57:22]
  reg  valid_6_7; // @[Cache.scala 57:22]
  reg  valid_7_0; // @[Cache.scala 57:22]
  reg  valid_7_1; // @[Cache.scala 57:22]
  reg  valid_7_2; // @[Cache.scala 57:22]
  reg  valid_7_3; // @[Cache.scala 57:22]
  reg  valid_7_4; // @[Cache.scala 57:22]
  reg  valid_7_5; // @[Cache.scala 57:22]
  reg  valid_7_6; // @[Cache.scala 57:22]
  reg  valid_7_7; // @[Cache.scala 57:22]
  reg  dirty_0_0; // @[Cache.scala 58:22]
  reg  dirty_0_1; // @[Cache.scala 58:22]
  reg  dirty_0_2; // @[Cache.scala 58:22]
  reg  dirty_0_3; // @[Cache.scala 58:22]
  reg  dirty_0_4; // @[Cache.scala 58:22]
  reg  dirty_0_5; // @[Cache.scala 58:22]
  reg  dirty_0_6; // @[Cache.scala 58:22]
  reg  dirty_0_7; // @[Cache.scala 58:22]
  reg  dirty_1_0; // @[Cache.scala 58:22]
  reg  dirty_1_1; // @[Cache.scala 58:22]
  reg  dirty_1_2; // @[Cache.scala 58:22]
  reg  dirty_1_3; // @[Cache.scala 58:22]
  reg  dirty_1_4; // @[Cache.scala 58:22]
  reg  dirty_1_5; // @[Cache.scala 58:22]
  reg  dirty_1_6; // @[Cache.scala 58:22]
  reg  dirty_1_7; // @[Cache.scala 58:22]
  reg  dirty_2_0; // @[Cache.scala 58:22]
  reg  dirty_2_1; // @[Cache.scala 58:22]
  reg  dirty_2_2; // @[Cache.scala 58:22]
  reg  dirty_2_3; // @[Cache.scala 58:22]
  reg  dirty_2_4; // @[Cache.scala 58:22]
  reg  dirty_2_5; // @[Cache.scala 58:22]
  reg  dirty_2_6; // @[Cache.scala 58:22]
  reg  dirty_2_7; // @[Cache.scala 58:22]
  reg  dirty_3_0; // @[Cache.scala 58:22]
  reg  dirty_3_1; // @[Cache.scala 58:22]
  reg  dirty_3_2; // @[Cache.scala 58:22]
  reg  dirty_3_3; // @[Cache.scala 58:22]
  reg  dirty_3_4; // @[Cache.scala 58:22]
  reg  dirty_3_5; // @[Cache.scala 58:22]
  reg  dirty_3_6; // @[Cache.scala 58:22]
  reg  dirty_3_7; // @[Cache.scala 58:22]
  reg  dirty_4_0; // @[Cache.scala 58:22]
  reg  dirty_4_1; // @[Cache.scala 58:22]
  reg  dirty_4_2; // @[Cache.scala 58:22]
  reg  dirty_4_3; // @[Cache.scala 58:22]
  reg  dirty_4_4; // @[Cache.scala 58:22]
  reg  dirty_4_5; // @[Cache.scala 58:22]
  reg  dirty_4_6; // @[Cache.scala 58:22]
  reg  dirty_4_7; // @[Cache.scala 58:22]
  reg  dirty_5_0; // @[Cache.scala 58:22]
  reg  dirty_5_1; // @[Cache.scala 58:22]
  reg  dirty_5_2; // @[Cache.scala 58:22]
  reg  dirty_5_3; // @[Cache.scala 58:22]
  reg  dirty_5_4; // @[Cache.scala 58:22]
  reg  dirty_5_5; // @[Cache.scala 58:22]
  reg  dirty_5_6; // @[Cache.scala 58:22]
  reg  dirty_5_7; // @[Cache.scala 58:22]
  reg  dirty_6_0; // @[Cache.scala 58:22]
  reg  dirty_6_1; // @[Cache.scala 58:22]
  reg  dirty_6_2; // @[Cache.scala 58:22]
  reg  dirty_6_3; // @[Cache.scala 58:22]
  reg  dirty_6_4; // @[Cache.scala 58:22]
  reg  dirty_6_5; // @[Cache.scala 58:22]
  reg  dirty_6_6; // @[Cache.scala 58:22]
  reg  dirty_6_7; // @[Cache.scala 58:22]
  reg  dirty_7_0; // @[Cache.scala 58:22]
  reg  dirty_7_1; // @[Cache.scala 58:22]
  reg  dirty_7_2; // @[Cache.scala 58:22]
  reg  dirty_7_3; // @[Cache.scala 58:22]
  reg  dirty_7_4; // @[Cache.scala 58:22]
  reg  dirty_7_5; // @[Cache.scala 58:22]
  reg  dirty_7_6; // @[Cache.scala 58:22]
  reg  dirty_7_7; // @[Cache.scala 58:22]
  wire [2:0] line_addr = io_addr[4:2]; // @[Cache.scala 64:26]
  wire [2:0] set_addr = io_addr[7:5]; // @[Cache.scala 65:25]
  wire [5:0] tag_addr = io_addr[13:8]; // @[Cache.scala 66:25]
  reg [2:0] mem_rd_set_addr; // @[Cache.scala 70:32]
  reg [5:0] mem_rd_tag_addr; // @[Cache.scala 71:32]
  wire [8:0] mem_rd_addr = {mem_rd_tag_addr,mem_rd_set_addr}; // @[Cat.scala 31:58]
  reg [8:0] mem_wr_addr; // @[Cache.scala 73:28]
  wire  _T = io_w_req | io_r_req; // @[Cache.scala 84:17]
  wire  _GEN_1 = 3'h1 == set_addr ? valid_1_0 : valid_0_0; // @[Cache.scala 88:{32,32}]
  wire  _GEN_2 = 3'h2 == set_addr ? valid_2_0 : _GEN_1; // @[Cache.scala 88:{32,32}]
  wire  _GEN_3 = 3'h3 == set_addr ? valid_3_0 : _GEN_2; // @[Cache.scala 88:{32,32}]
  wire  _GEN_4 = 3'h4 == set_addr ? valid_4_0 : _GEN_3; // @[Cache.scala 88:{32,32}]
  wire  _GEN_5 = 3'h5 == set_addr ? valid_5_0 : _GEN_4; // @[Cache.scala 88:{32,32}]
  wire  _GEN_6 = 3'h6 == set_addr ? valid_6_0 : _GEN_5; // @[Cache.scala 88:{32,32}]
  wire  _GEN_7 = 3'h7 == set_addr ? valid_7_0 : _GEN_6; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_9 = 3'h1 == set_addr ? cache_tags_1_0 : cache_tags_0_0; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_10 = 3'h2 == set_addr ? cache_tags_2_0 : _GEN_9; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_11 = 3'h3 == set_addr ? cache_tags_3_0 : _GEN_10; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_12 = 3'h4 == set_addr ? cache_tags_4_0 : _GEN_11; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_13 = 3'h5 == set_addr ? cache_tags_5_0 : _GEN_12; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_14 = 3'h6 == set_addr ? cache_tags_6_0 : _GEN_13; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_15 = 3'h7 == set_addr ? cache_tags_7_0 : _GEN_14; // @[Cache.scala 88:{70,70}]
  wire  _GEN_19 = 3'h1 == set_addr ? valid_1_1 : valid_0_1; // @[Cache.scala 88:{32,32}]
  wire  _GEN_20 = 3'h2 == set_addr ? valid_2_1 : _GEN_19; // @[Cache.scala 88:{32,32}]
  wire  _GEN_21 = 3'h3 == set_addr ? valid_3_1 : _GEN_20; // @[Cache.scala 88:{32,32}]
  wire  _GEN_22 = 3'h4 == set_addr ? valid_4_1 : _GEN_21; // @[Cache.scala 88:{32,32}]
  wire  _GEN_23 = 3'h5 == set_addr ? valid_5_1 : _GEN_22; // @[Cache.scala 88:{32,32}]
  wire  _GEN_24 = 3'h6 == set_addr ? valid_6_1 : _GEN_23; // @[Cache.scala 88:{32,32}]
  wire  _GEN_25 = 3'h7 == set_addr ? valid_7_1 : _GEN_24; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_27 = 3'h1 == set_addr ? cache_tags_1_1 : cache_tags_0_1; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_28 = 3'h2 == set_addr ? cache_tags_2_1 : _GEN_27; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_29 = 3'h3 == set_addr ? cache_tags_3_1 : _GEN_28; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_30 = 3'h4 == set_addr ? cache_tags_4_1 : _GEN_29; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_31 = 3'h5 == set_addr ? cache_tags_5_1 : _GEN_30; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_32 = 3'h6 == set_addr ? cache_tags_6_1 : _GEN_31; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_33 = 3'h7 == set_addr ? cache_tags_7_1 : _GEN_32; // @[Cache.scala 88:{70,70}]
  wire  _T_6 = _GEN_25 & _GEN_33 == tag_addr; // @[Cache.scala 88:42]
  wire  _GEN_37 = 3'h1 == set_addr ? valid_1_2 : valid_0_2; // @[Cache.scala 88:{32,32}]
  wire  _GEN_38 = 3'h2 == set_addr ? valid_2_2 : _GEN_37; // @[Cache.scala 88:{32,32}]
  wire  _GEN_39 = 3'h3 == set_addr ? valid_3_2 : _GEN_38; // @[Cache.scala 88:{32,32}]
  wire  _GEN_40 = 3'h4 == set_addr ? valid_4_2 : _GEN_39; // @[Cache.scala 88:{32,32}]
  wire  _GEN_41 = 3'h5 == set_addr ? valid_5_2 : _GEN_40; // @[Cache.scala 88:{32,32}]
  wire  _GEN_42 = 3'h6 == set_addr ? valid_6_2 : _GEN_41; // @[Cache.scala 88:{32,32}]
  wire  _GEN_43 = 3'h7 == set_addr ? valid_7_2 : _GEN_42; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_45 = 3'h1 == set_addr ? cache_tags_1_2 : cache_tags_0_2; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_46 = 3'h2 == set_addr ? cache_tags_2_2 : _GEN_45; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_47 = 3'h3 == set_addr ? cache_tags_3_2 : _GEN_46; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_48 = 3'h4 == set_addr ? cache_tags_4_2 : _GEN_47; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_49 = 3'h5 == set_addr ? cache_tags_5_2 : _GEN_48; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_50 = 3'h6 == set_addr ? cache_tags_6_2 : _GEN_49; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_51 = 3'h7 == set_addr ? cache_tags_7_2 : _GEN_50; // @[Cache.scala 88:{70,70}]
  wire [1:0] _GEN_53 = _GEN_43 & _GEN_51 == tag_addr ? 2'h2 : {{1'd0}, _T_6}; // @[Cache.scala 88:82 90:17]
  wire  _GEN_55 = 3'h1 == set_addr ? valid_1_3 : valid_0_3; // @[Cache.scala 88:{32,32}]
  wire  _GEN_56 = 3'h2 == set_addr ? valid_2_3 : _GEN_55; // @[Cache.scala 88:{32,32}]
  wire  _GEN_57 = 3'h3 == set_addr ? valid_3_3 : _GEN_56; // @[Cache.scala 88:{32,32}]
  wire  _GEN_58 = 3'h4 == set_addr ? valid_4_3 : _GEN_57; // @[Cache.scala 88:{32,32}]
  wire  _GEN_59 = 3'h5 == set_addr ? valid_5_3 : _GEN_58; // @[Cache.scala 88:{32,32}]
  wire  _GEN_60 = 3'h6 == set_addr ? valid_6_3 : _GEN_59; // @[Cache.scala 88:{32,32}]
  wire  _GEN_61 = 3'h7 == set_addr ? valid_7_3 : _GEN_60; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_63 = 3'h1 == set_addr ? cache_tags_1_3 : cache_tags_0_3; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_64 = 3'h2 == set_addr ? cache_tags_2_3 : _GEN_63; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_65 = 3'h3 == set_addr ? cache_tags_3_3 : _GEN_64; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_66 = 3'h4 == set_addr ? cache_tags_4_3 : _GEN_65; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_67 = 3'h5 == set_addr ? cache_tags_5_3 : _GEN_66; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_68 = 3'h6 == set_addr ? cache_tags_6_3 : _GEN_67; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_69 = 3'h7 == set_addr ? cache_tags_7_3 : _GEN_68; // @[Cache.scala 88:{70,70}]
  wire [1:0] _GEN_71 = _GEN_61 & _GEN_69 == tag_addr ? 2'h3 : _GEN_53; // @[Cache.scala 88:82 90:17]
  wire  _GEN_73 = 3'h1 == set_addr ? valid_1_4 : valid_0_4; // @[Cache.scala 88:{32,32}]
  wire  _GEN_74 = 3'h2 == set_addr ? valid_2_4 : _GEN_73; // @[Cache.scala 88:{32,32}]
  wire  _GEN_75 = 3'h3 == set_addr ? valid_3_4 : _GEN_74; // @[Cache.scala 88:{32,32}]
  wire  _GEN_76 = 3'h4 == set_addr ? valid_4_4 : _GEN_75; // @[Cache.scala 88:{32,32}]
  wire  _GEN_77 = 3'h5 == set_addr ? valid_5_4 : _GEN_76; // @[Cache.scala 88:{32,32}]
  wire  _GEN_78 = 3'h6 == set_addr ? valid_6_4 : _GEN_77; // @[Cache.scala 88:{32,32}]
  wire  _GEN_79 = 3'h7 == set_addr ? valid_7_4 : _GEN_78; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_81 = 3'h1 == set_addr ? cache_tags_1_4 : cache_tags_0_4; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_82 = 3'h2 == set_addr ? cache_tags_2_4 : _GEN_81; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_83 = 3'h3 == set_addr ? cache_tags_3_4 : _GEN_82; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_84 = 3'h4 == set_addr ? cache_tags_4_4 : _GEN_83; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_85 = 3'h5 == set_addr ? cache_tags_5_4 : _GEN_84; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_86 = 3'h6 == set_addr ? cache_tags_6_4 : _GEN_85; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_87 = 3'h7 == set_addr ? cache_tags_7_4 : _GEN_86; // @[Cache.scala 88:{70,70}]
  wire [2:0] _GEN_89 = _GEN_79 & _GEN_87 == tag_addr ? 3'h4 : {{1'd0}, _GEN_71}; // @[Cache.scala 88:82 90:17]
  wire  _GEN_91 = 3'h1 == set_addr ? valid_1_5 : valid_0_5; // @[Cache.scala 88:{32,32}]
  wire  _GEN_92 = 3'h2 == set_addr ? valid_2_5 : _GEN_91; // @[Cache.scala 88:{32,32}]
  wire  _GEN_93 = 3'h3 == set_addr ? valid_3_5 : _GEN_92; // @[Cache.scala 88:{32,32}]
  wire  _GEN_94 = 3'h4 == set_addr ? valid_4_5 : _GEN_93; // @[Cache.scala 88:{32,32}]
  wire  _GEN_95 = 3'h5 == set_addr ? valid_5_5 : _GEN_94; // @[Cache.scala 88:{32,32}]
  wire  _GEN_96 = 3'h6 == set_addr ? valid_6_5 : _GEN_95; // @[Cache.scala 88:{32,32}]
  wire  _GEN_97 = 3'h7 == set_addr ? valid_7_5 : _GEN_96; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_99 = 3'h1 == set_addr ? cache_tags_1_5 : cache_tags_0_5; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_100 = 3'h2 == set_addr ? cache_tags_2_5 : _GEN_99; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_101 = 3'h3 == set_addr ? cache_tags_3_5 : _GEN_100; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_102 = 3'h4 == set_addr ? cache_tags_4_5 : _GEN_101; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_103 = 3'h5 == set_addr ? cache_tags_5_5 : _GEN_102; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_104 = 3'h6 == set_addr ? cache_tags_6_5 : _GEN_103; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_105 = 3'h7 == set_addr ? cache_tags_7_5 : _GEN_104; // @[Cache.scala 88:{70,70}]
  wire [2:0] _GEN_107 = _GEN_97 & _GEN_105 == tag_addr ? 3'h5 : _GEN_89; // @[Cache.scala 88:82 90:17]
  wire  _GEN_109 = 3'h1 == set_addr ? valid_1_6 : valid_0_6; // @[Cache.scala 88:{32,32}]
  wire  _GEN_110 = 3'h2 == set_addr ? valid_2_6 : _GEN_109; // @[Cache.scala 88:{32,32}]
  wire  _GEN_111 = 3'h3 == set_addr ? valid_3_6 : _GEN_110; // @[Cache.scala 88:{32,32}]
  wire  _GEN_112 = 3'h4 == set_addr ? valid_4_6 : _GEN_111; // @[Cache.scala 88:{32,32}]
  wire  _GEN_113 = 3'h5 == set_addr ? valid_5_6 : _GEN_112; // @[Cache.scala 88:{32,32}]
  wire  _GEN_114 = 3'h6 == set_addr ? valid_6_6 : _GEN_113; // @[Cache.scala 88:{32,32}]
  wire  _GEN_115 = 3'h7 == set_addr ? valid_7_6 : _GEN_114; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_117 = 3'h1 == set_addr ? cache_tags_1_6 : cache_tags_0_6; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_118 = 3'h2 == set_addr ? cache_tags_2_6 : _GEN_117; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_119 = 3'h3 == set_addr ? cache_tags_3_6 : _GEN_118; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_120 = 3'h4 == set_addr ? cache_tags_4_6 : _GEN_119; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_121 = 3'h5 == set_addr ? cache_tags_5_6 : _GEN_120; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_122 = 3'h6 == set_addr ? cache_tags_6_6 : _GEN_121; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_123 = 3'h7 == set_addr ? cache_tags_7_6 : _GEN_122; // @[Cache.scala 88:{70,70}]
  wire [2:0] _GEN_125 = _GEN_115 & _GEN_123 == tag_addr ? 3'h6 : _GEN_107; // @[Cache.scala 88:82 90:17]
  wire  _GEN_127 = 3'h1 == set_addr ? valid_1_7 : valid_0_7; // @[Cache.scala 88:{32,32}]
  wire  _GEN_128 = 3'h2 == set_addr ? valid_2_7 : _GEN_127; // @[Cache.scala 88:{32,32}]
  wire  _GEN_129 = 3'h3 == set_addr ? valid_3_7 : _GEN_128; // @[Cache.scala 88:{32,32}]
  wire  _GEN_130 = 3'h4 == set_addr ? valid_4_7 : _GEN_129; // @[Cache.scala 88:{32,32}]
  wire  _GEN_131 = 3'h5 == set_addr ? valid_5_7 : _GEN_130; // @[Cache.scala 88:{32,32}]
  wire  _GEN_132 = 3'h6 == set_addr ? valid_6_7 : _GEN_131; // @[Cache.scala 88:{32,32}]
  wire  _GEN_133 = 3'h7 == set_addr ? valid_7_7 : _GEN_132; // @[Cache.scala 88:{32,32}]
  wire [5:0] _GEN_135 = 3'h1 == set_addr ? cache_tags_1_7 : cache_tags_0_7; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_136 = 3'h2 == set_addr ? cache_tags_2_7 : _GEN_135; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_137 = 3'h3 == set_addr ? cache_tags_3_7 : _GEN_136; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_138 = 3'h4 == set_addr ? cache_tags_4_7 : _GEN_137; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_139 = 3'h5 == set_addr ? cache_tags_5_7 : _GEN_138; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_140 = 3'h6 == set_addr ? cache_tags_6_7 : _GEN_139; // @[Cache.scala 88:{70,70}]
  wire [5:0] _GEN_141 = 3'h7 == set_addr ? cache_tags_7_7 : _GEN_140; // @[Cache.scala 88:{70,70}]
  wire  _GEN_142 = _GEN_133 & _GEN_141 == tag_addr | (_GEN_115 & _GEN_123 == tag_addr | (_GEN_97 & _GEN_105 == tag_addr
     | (_GEN_79 & _GEN_87 == tag_addr | (_GEN_61 & _GEN_69 == tag_addr | (_GEN_43 & _GEN_51 == tag_addr | (_GEN_25 &
    _GEN_33 == tag_addr | _GEN_7 & _GEN_15 == tag_addr)))))); // @[Cache.scala 88:82 89:19]
  wire [2:0] _GEN_143 = _GEN_133 & _GEN_141 == tag_addr ? 3'h7 : _GEN_125; // @[Cache.scala 88:82 90:17]
  wire  cache_Hit = (io_w_req | io_r_req) & _GEN_142; // @[Cache.scala 84:28]
  wire [2:0] way_hit = io_w_req | io_r_req ? _GEN_143 : 3'h0; // @[Cache.scala 84:28]
  reg [1:0] cacheState; // @[Cache.scala 96:27]
  reg [31:0] FIFO_Choice_0; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_1; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_2; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_3; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_4; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_5; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_6; // @[Cache.scala 103:30]
  reg [31:0] FIFO_Choice_7; // @[Cache.scala 103:30]
  wire  _T_27 = 2'h0 == cacheState; // @[Cache.scala 104:23]
  wire [31:0] _GEN_147 = 3'h1 == set_addr ? FIFO_Choice_1 : FIFO_Choice_0; // @[Cache.scala 106:{23,23}]
  wire [31:0] _GEN_148 = 3'h2 == set_addr ? FIFO_Choice_2 : _GEN_147; // @[Cache.scala 106:{23,23}]
  wire [31:0] _GEN_149 = 3'h3 == set_addr ? FIFO_Choice_3 : _GEN_148; // @[Cache.scala 106:{23,23}]
  wire [31:0] _GEN_150 = 3'h4 == set_addr ? FIFO_Choice_4 : _GEN_149; // @[Cache.scala 106:{23,23}]
  wire [31:0] _GEN_151 = 3'h5 == set_addr ? FIFO_Choice_5 : _GEN_150; // @[Cache.scala 106:{23,23}]
  wire [31:0] _GEN_152 = 3'h6 == set_addr ? FIFO_Choice_6 : _GEN_151; // @[Cache.scala 106:{23,23}]
  wire [31:0] _GEN_153 = 3'h7 == set_addr ? FIFO_Choice_7 : _GEN_152; // @[Cache.scala 106:{23,23}]
  wire  _T_30 = 2'h3 == cacheState; // @[Cache.scala 104:23]
  wire [31:0] _FIFO_Choice_T_1 = _GEN_153 + 32'h1; // @[Cache.scala 109:57]
  wire [31:0] _GEN_0 = _FIFO_Choice_T_1 % 32'h8; // @[Cache.scala 109:63]
  wire [31:0] _FIFO_Choice_set_addr_1 = {{28'd0}, _GEN_0[3:0]}; // @[Cache.scala 109:{31,31}]
  wire [31:0] _GEN_170 = 2'h0 == cacheState ? _GEN_153 : 32'h0; // @[Cache.scala 104:23 106:23]
  reg [31:0] mem_wr_line_0; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_1; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_2; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_3; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_4; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_5; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_6; // @[Cache.scala 124:28]
  reg [31:0] mem_wr_line_7; // @[Cache.scala 124:28]
  wire  _GEN_9835 = 3'h0 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9837 = 3'h0 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9838 = 3'h1 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_180 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_0_0_1 : CacheMem_0_0_0; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9842 = 3'h2 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_181 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_0_0_2 : _GEN_180; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9846 = 3'h3 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_182 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_0_0_3 : _GEN_181; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9850 = 3'h4 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_183 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_0_0_4 : _GEN_182; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9854 = 3'h5 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_184 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_0_0_5 : _GEN_183; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9858 = 3'h6 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_185 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_0_0_6 : _GEN_184; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9862 = 3'h7 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_186 = 3'h0 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_0_0_7 : _GEN_185; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9865 = 3'h0 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9866 = 3'h0 == line_addr; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_187 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_0_1_0 : _GEN_186; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_188 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_0_1_1 : _GEN_187; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_189 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_0_1_2 : _GEN_188; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_190 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_0_1_3 : _GEN_189; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_191 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_0_1_4 : _GEN_190; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_192 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_0_1_5 : _GEN_191; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_193 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_0_1_6 : _GEN_192; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_194 = 3'h0 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_0_1_7 : _GEN_193; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9897 = 3'h0 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_195 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_0_2_0 : _GEN_194; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_196 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_0_2_1 : _GEN_195; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_197 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_0_2_2 : _GEN_196; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_198 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_0_2_3 : _GEN_197; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_199 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_0_2_4 : _GEN_198; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_200 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_0_2_5 : _GEN_199; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_201 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_0_2_6 : _GEN_200; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_202 = 3'h0 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_0_2_7 : _GEN_201; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9929 = 3'h0 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_203 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_0_3_0 : _GEN_202; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_204 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_0_3_1 : _GEN_203; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_205 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_0_3_2 : _GEN_204; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_206 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_0_3_3 : _GEN_205; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_207 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_0_3_4 : _GEN_206; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_208 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_0_3_5 : _GEN_207; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_209 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_0_3_6 : _GEN_208; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_210 = 3'h0 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_0_3_7 : _GEN_209; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9961 = 3'h0 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_211 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_0_4_0 : _GEN_210; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_212 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_0_4_1 : _GEN_211; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_213 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_0_4_2 : _GEN_212; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_214 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_0_4_3 : _GEN_213; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_215 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_0_4_4 : _GEN_214; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_216 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_0_4_5 : _GEN_215; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_217 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_0_4_6 : _GEN_216; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_218 = 3'h0 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_0_4_7 : _GEN_217; // @[Cache.scala 131:{15,15}]
  wire  _GEN_9993 = 3'h0 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_219 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_0_5_0 : _GEN_218; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_220 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_0_5_1 : _GEN_219; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_221 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_0_5_2 : _GEN_220; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_222 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_0_5_3 : _GEN_221; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_223 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_0_5_4 : _GEN_222; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_224 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_0_5_5 : _GEN_223; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_225 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_0_5_6 : _GEN_224; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_226 = 3'h0 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_0_5_7 : _GEN_225; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10025 = 3'h0 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_227 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_0_6_0 : _GEN_226; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_228 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_0_6_1 : _GEN_227; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_229 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_0_6_2 : _GEN_228; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_230 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_0_6_3 : _GEN_229; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_231 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_0_6_4 : _GEN_230; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_232 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_0_6_5 : _GEN_231; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_233 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_0_6_6 : _GEN_232; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_234 = 3'h0 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_0_6_7 : _GEN_233; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10057 = 3'h0 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_235 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_0_7_0 : _GEN_234; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_236 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_0_7_1 : _GEN_235; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_237 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_0_7_2 : _GEN_236; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_238 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_0_7_3 : _GEN_237; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_239 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_0_7_4 : _GEN_238; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_240 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_0_7_5 : _GEN_239; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_241 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_0_7_6 : _GEN_240; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_242 = 3'h0 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_0_7_7 : _GEN_241; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10087 = 3'h1 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10089 = 3'h1 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_243 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_1_0_0 : _GEN_242; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_244 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_1_0_1 : _GEN_243; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_245 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_1_0_2 : _GEN_244; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_246 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_1_0_3 : _GEN_245; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_247 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_1_0_4 : _GEN_246; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_248 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_1_0_5 : _GEN_247; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_249 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_1_0_6 : _GEN_248; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_250 = 3'h1 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_1_0_7 : _GEN_249; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10121 = 3'h1 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_251 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_1_1_0 : _GEN_250; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_252 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_1_1_1 : _GEN_251; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_253 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_1_1_2 : _GEN_252; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_254 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_1_1_3 : _GEN_253; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_255 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_1_1_4 : _GEN_254; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_256 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_1_1_5 : _GEN_255; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_257 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_1_1_6 : _GEN_256; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_258 = 3'h1 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_1_1_7 : _GEN_257; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10153 = 3'h1 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_259 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_1_2_0 : _GEN_258; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_260 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_1_2_1 : _GEN_259; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_261 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_1_2_2 : _GEN_260; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_262 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_1_2_3 : _GEN_261; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_263 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_1_2_4 : _GEN_262; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_264 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_1_2_5 : _GEN_263; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_265 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_1_2_6 : _GEN_264; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_266 = 3'h1 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_1_2_7 : _GEN_265; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10185 = 3'h1 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_267 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_1_3_0 : _GEN_266; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_268 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_1_3_1 : _GEN_267; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_269 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_1_3_2 : _GEN_268; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_270 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_1_3_3 : _GEN_269; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_271 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_1_3_4 : _GEN_270; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_272 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_1_3_5 : _GEN_271; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_273 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_1_3_6 : _GEN_272; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_274 = 3'h1 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_1_3_7 : _GEN_273; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10217 = 3'h1 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_275 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_1_4_0 : _GEN_274; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_276 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_1_4_1 : _GEN_275; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_277 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_1_4_2 : _GEN_276; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_278 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_1_4_3 : _GEN_277; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_279 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_1_4_4 : _GEN_278; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_280 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_1_4_5 : _GEN_279; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_281 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_1_4_6 : _GEN_280; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_282 = 3'h1 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_1_4_7 : _GEN_281; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10249 = 3'h1 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_283 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_1_5_0 : _GEN_282; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_284 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_1_5_1 : _GEN_283; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_285 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_1_5_2 : _GEN_284; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_286 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_1_5_3 : _GEN_285; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_287 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_1_5_4 : _GEN_286; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_288 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_1_5_5 : _GEN_287; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_289 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_1_5_6 : _GEN_288; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_290 = 3'h1 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_1_5_7 : _GEN_289; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10281 = 3'h1 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_291 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_1_6_0 : _GEN_290; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_292 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_1_6_1 : _GEN_291; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_293 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_1_6_2 : _GEN_292; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_294 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_1_6_3 : _GEN_293; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_295 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_1_6_4 : _GEN_294; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_296 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_1_6_5 : _GEN_295; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_297 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_1_6_6 : _GEN_296; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_298 = 3'h1 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_1_6_7 : _GEN_297; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10313 = 3'h1 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_299 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_1_7_0 : _GEN_298; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_300 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_1_7_1 : _GEN_299; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_301 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_1_7_2 : _GEN_300; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_302 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_1_7_3 : _GEN_301; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_303 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_1_7_4 : _GEN_302; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_304 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_1_7_5 : _GEN_303; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_305 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_1_7_6 : _GEN_304; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_306 = 3'h1 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_1_7_7 : _GEN_305; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10343 = 3'h2 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10345 = 3'h2 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_307 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_2_0_0 : _GEN_306; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_308 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_2_0_1 : _GEN_307; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_309 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_2_0_2 : _GEN_308; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_310 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_2_0_3 : _GEN_309; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_311 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_2_0_4 : _GEN_310; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_312 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_2_0_5 : _GEN_311; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_313 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_2_0_6 : _GEN_312; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_314 = 3'h2 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_2_0_7 : _GEN_313; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10377 = 3'h2 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_315 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_2_1_0 : _GEN_314; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_316 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_2_1_1 : _GEN_315; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_317 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_2_1_2 : _GEN_316; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_318 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_2_1_3 : _GEN_317; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_319 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_2_1_4 : _GEN_318; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_320 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_2_1_5 : _GEN_319; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_321 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_2_1_6 : _GEN_320; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_322 = 3'h2 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_2_1_7 : _GEN_321; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10409 = 3'h2 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_323 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_2_2_0 : _GEN_322; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_324 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_2_2_1 : _GEN_323; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_325 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_2_2_2 : _GEN_324; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_326 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_2_2_3 : _GEN_325; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_327 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_2_2_4 : _GEN_326; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_328 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_2_2_5 : _GEN_327; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_329 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_2_2_6 : _GEN_328; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_330 = 3'h2 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_2_2_7 : _GEN_329; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10441 = 3'h2 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_331 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_2_3_0 : _GEN_330; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_332 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_2_3_1 : _GEN_331; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_333 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_2_3_2 : _GEN_332; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_334 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_2_3_3 : _GEN_333; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_335 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_2_3_4 : _GEN_334; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_336 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_2_3_5 : _GEN_335; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_337 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_2_3_6 : _GEN_336; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_338 = 3'h2 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_2_3_7 : _GEN_337; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10473 = 3'h2 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_339 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_2_4_0 : _GEN_338; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_340 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_2_4_1 : _GEN_339; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_341 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_2_4_2 : _GEN_340; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_342 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_2_4_3 : _GEN_341; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_343 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_2_4_4 : _GEN_342; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_344 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_2_4_5 : _GEN_343; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_345 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_2_4_6 : _GEN_344; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_346 = 3'h2 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_2_4_7 : _GEN_345; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10505 = 3'h2 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_347 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_2_5_0 : _GEN_346; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_348 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_2_5_1 : _GEN_347; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_349 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_2_5_2 : _GEN_348; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_350 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_2_5_3 : _GEN_349; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_351 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_2_5_4 : _GEN_350; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_352 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_2_5_5 : _GEN_351; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_353 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_2_5_6 : _GEN_352; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_354 = 3'h2 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_2_5_7 : _GEN_353; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10537 = 3'h2 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_355 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_2_6_0 : _GEN_354; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_356 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_2_6_1 : _GEN_355; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_357 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_2_6_2 : _GEN_356; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_358 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_2_6_3 : _GEN_357; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_359 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_2_6_4 : _GEN_358; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_360 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_2_6_5 : _GEN_359; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_361 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_2_6_6 : _GEN_360; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_362 = 3'h2 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_2_6_7 : _GEN_361; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10569 = 3'h2 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_363 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_2_7_0 : _GEN_362; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_364 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_2_7_1 : _GEN_363; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_365 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_2_7_2 : _GEN_364; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_366 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_2_7_3 : _GEN_365; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_367 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_2_7_4 : _GEN_366; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_368 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_2_7_5 : _GEN_367; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_369 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_2_7_6 : _GEN_368; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_370 = 3'h2 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_2_7_7 : _GEN_369; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10599 = 3'h3 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10601 = 3'h3 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_371 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_3_0_0 : _GEN_370; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_372 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_3_0_1 : _GEN_371; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_373 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_3_0_2 : _GEN_372; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_374 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_3_0_3 : _GEN_373; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_375 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_3_0_4 : _GEN_374; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_376 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_3_0_5 : _GEN_375; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_377 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_3_0_6 : _GEN_376; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_378 = 3'h3 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_3_0_7 : _GEN_377; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10633 = 3'h3 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_379 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_3_1_0 : _GEN_378; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_380 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_3_1_1 : _GEN_379; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_381 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_3_1_2 : _GEN_380; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_382 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_3_1_3 : _GEN_381; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_383 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_3_1_4 : _GEN_382; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_384 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_3_1_5 : _GEN_383; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_385 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_3_1_6 : _GEN_384; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_386 = 3'h3 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_3_1_7 : _GEN_385; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10665 = 3'h3 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_387 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_3_2_0 : _GEN_386; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_388 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_3_2_1 : _GEN_387; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_389 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_3_2_2 : _GEN_388; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_390 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_3_2_3 : _GEN_389; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_391 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_3_2_4 : _GEN_390; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_392 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_3_2_5 : _GEN_391; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_393 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_3_2_6 : _GEN_392; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_394 = 3'h3 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_3_2_7 : _GEN_393; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10697 = 3'h3 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_395 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_3_3_0 : _GEN_394; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_396 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_3_3_1 : _GEN_395; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_397 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_3_3_2 : _GEN_396; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_398 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_3_3_3 : _GEN_397; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_399 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_3_3_4 : _GEN_398; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_400 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_3_3_5 : _GEN_399; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_401 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_3_3_6 : _GEN_400; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_402 = 3'h3 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_3_3_7 : _GEN_401; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10729 = 3'h3 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_403 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_3_4_0 : _GEN_402; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_404 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_3_4_1 : _GEN_403; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_405 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_3_4_2 : _GEN_404; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_406 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_3_4_3 : _GEN_405; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_407 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_3_4_4 : _GEN_406; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_408 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_3_4_5 : _GEN_407; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_409 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_3_4_6 : _GEN_408; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_410 = 3'h3 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_3_4_7 : _GEN_409; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10761 = 3'h3 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_411 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_3_5_0 : _GEN_410; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_412 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_3_5_1 : _GEN_411; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_413 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_3_5_2 : _GEN_412; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_414 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_3_5_3 : _GEN_413; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_415 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_3_5_4 : _GEN_414; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_416 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_3_5_5 : _GEN_415; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_417 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_3_5_6 : _GEN_416; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_418 = 3'h3 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_3_5_7 : _GEN_417; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10793 = 3'h3 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_419 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_3_6_0 : _GEN_418; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_420 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_3_6_1 : _GEN_419; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_421 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_3_6_2 : _GEN_420; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_422 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_3_6_3 : _GEN_421; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_423 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_3_6_4 : _GEN_422; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_424 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_3_6_5 : _GEN_423; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_425 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_3_6_6 : _GEN_424; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_426 = 3'h3 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_3_6_7 : _GEN_425; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10825 = 3'h3 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_427 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_3_7_0 : _GEN_426; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_428 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_3_7_1 : _GEN_427; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_429 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_3_7_2 : _GEN_428; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_430 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_3_7_3 : _GEN_429; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_431 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_3_7_4 : _GEN_430; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_432 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_3_7_5 : _GEN_431; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_433 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_3_7_6 : _GEN_432; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_434 = 3'h3 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_3_7_7 : _GEN_433; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10855 = 3'h4 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10857 = 3'h4 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_435 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_4_0_0 : _GEN_434; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_436 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_4_0_1 : _GEN_435; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_437 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_4_0_2 : _GEN_436; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_438 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_4_0_3 : _GEN_437; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_439 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_4_0_4 : _GEN_438; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_440 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_4_0_5 : _GEN_439; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_441 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_4_0_6 : _GEN_440; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_442 = 3'h4 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_4_0_7 : _GEN_441; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10889 = 3'h4 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_443 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_4_1_0 : _GEN_442; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_444 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_4_1_1 : _GEN_443; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_445 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_4_1_2 : _GEN_444; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_446 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_4_1_3 : _GEN_445; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_447 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_4_1_4 : _GEN_446; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_448 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_4_1_5 : _GEN_447; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_449 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_4_1_6 : _GEN_448; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_450 = 3'h4 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_4_1_7 : _GEN_449; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10921 = 3'h4 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_451 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_4_2_0 : _GEN_450; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_452 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_4_2_1 : _GEN_451; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_453 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_4_2_2 : _GEN_452; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_454 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_4_2_3 : _GEN_453; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_455 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_4_2_4 : _GEN_454; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_456 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_4_2_5 : _GEN_455; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_457 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_4_2_6 : _GEN_456; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_458 = 3'h4 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_4_2_7 : _GEN_457; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10953 = 3'h4 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_459 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_4_3_0 : _GEN_458; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_460 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_4_3_1 : _GEN_459; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_461 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_4_3_2 : _GEN_460; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_462 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_4_3_3 : _GEN_461; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_463 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_4_3_4 : _GEN_462; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_464 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_4_3_5 : _GEN_463; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_465 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_4_3_6 : _GEN_464; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_466 = 3'h4 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_4_3_7 : _GEN_465; // @[Cache.scala 131:{15,15}]
  wire  _GEN_10985 = 3'h4 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_467 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_4_4_0 : _GEN_466; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_468 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_4_4_1 : _GEN_467; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_469 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_4_4_2 : _GEN_468; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_470 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_4_4_3 : _GEN_469; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_471 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_4_4_4 : _GEN_470; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_472 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_4_4_5 : _GEN_471; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_473 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_4_4_6 : _GEN_472; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_474 = 3'h4 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_4_4_7 : _GEN_473; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11017 = 3'h4 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_475 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_4_5_0 : _GEN_474; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_476 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_4_5_1 : _GEN_475; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_477 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_4_5_2 : _GEN_476; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_478 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_4_5_3 : _GEN_477; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_479 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_4_5_4 : _GEN_478; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_480 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_4_5_5 : _GEN_479; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_481 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_4_5_6 : _GEN_480; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_482 = 3'h4 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_4_5_7 : _GEN_481; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11049 = 3'h4 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_483 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_4_6_0 : _GEN_482; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_484 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_4_6_1 : _GEN_483; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_485 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_4_6_2 : _GEN_484; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_486 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_4_6_3 : _GEN_485; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_487 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_4_6_4 : _GEN_486; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_488 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_4_6_5 : _GEN_487; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_489 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_4_6_6 : _GEN_488; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_490 = 3'h4 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_4_6_7 : _GEN_489; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11081 = 3'h4 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_491 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_4_7_0 : _GEN_490; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_492 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_4_7_1 : _GEN_491; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_493 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_4_7_2 : _GEN_492; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_494 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_4_7_3 : _GEN_493; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_495 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_4_7_4 : _GEN_494; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_496 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_4_7_5 : _GEN_495; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_497 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_4_7_6 : _GEN_496; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_498 = 3'h4 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_4_7_7 : _GEN_497; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11111 = 3'h5 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11113 = 3'h5 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_499 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_5_0_0 : _GEN_498; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_500 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_5_0_1 : _GEN_499; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_501 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_5_0_2 : _GEN_500; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_502 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_5_0_3 : _GEN_501; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_503 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_5_0_4 : _GEN_502; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_504 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_5_0_5 : _GEN_503; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_505 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_5_0_6 : _GEN_504; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_506 = 3'h5 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_5_0_7 : _GEN_505; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11145 = 3'h5 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_507 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_5_1_0 : _GEN_506; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_508 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_5_1_1 : _GEN_507; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_509 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_5_1_2 : _GEN_508; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_510 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_5_1_3 : _GEN_509; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_511 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_5_1_4 : _GEN_510; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_512 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_5_1_5 : _GEN_511; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_513 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_5_1_6 : _GEN_512; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_514 = 3'h5 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_5_1_7 : _GEN_513; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11177 = 3'h5 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_515 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_5_2_0 : _GEN_514; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_516 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_5_2_1 : _GEN_515; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_517 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_5_2_2 : _GEN_516; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_518 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_5_2_3 : _GEN_517; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_519 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_5_2_4 : _GEN_518; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_520 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_5_2_5 : _GEN_519; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_521 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_5_2_6 : _GEN_520; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_522 = 3'h5 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_5_2_7 : _GEN_521; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11209 = 3'h5 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_523 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_5_3_0 : _GEN_522; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_524 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_5_3_1 : _GEN_523; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_525 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_5_3_2 : _GEN_524; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_526 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_5_3_3 : _GEN_525; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_527 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_5_3_4 : _GEN_526; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_528 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_5_3_5 : _GEN_527; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_529 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_5_3_6 : _GEN_528; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_530 = 3'h5 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_5_3_7 : _GEN_529; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11241 = 3'h5 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_531 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_5_4_0 : _GEN_530; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_532 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_5_4_1 : _GEN_531; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_533 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_5_4_2 : _GEN_532; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_534 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_5_4_3 : _GEN_533; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_535 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_5_4_4 : _GEN_534; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_536 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_5_4_5 : _GEN_535; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_537 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_5_4_6 : _GEN_536; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_538 = 3'h5 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_5_4_7 : _GEN_537; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11273 = 3'h5 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_539 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_5_5_0 : _GEN_538; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_540 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_5_5_1 : _GEN_539; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_541 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_5_5_2 : _GEN_540; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_542 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_5_5_3 : _GEN_541; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_543 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_5_5_4 : _GEN_542; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_544 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_5_5_5 : _GEN_543; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_545 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_5_5_6 : _GEN_544; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_546 = 3'h5 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_5_5_7 : _GEN_545; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11305 = 3'h5 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_547 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_5_6_0 : _GEN_546; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_548 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_5_6_1 : _GEN_547; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_549 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_5_6_2 : _GEN_548; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_550 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_5_6_3 : _GEN_549; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_551 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_5_6_4 : _GEN_550; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_552 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_5_6_5 : _GEN_551; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_553 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_5_6_6 : _GEN_552; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_554 = 3'h5 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_5_6_7 : _GEN_553; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11337 = 3'h5 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_555 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_5_7_0 : _GEN_554; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_556 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_5_7_1 : _GEN_555; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_557 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_5_7_2 : _GEN_556; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_558 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_5_7_3 : _GEN_557; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_559 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_5_7_4 : _GEN_558; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_560 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_5_7_5 : _GEN_559; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_561 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_5_7_6 : _GEN_560; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_562 = 3'h5 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_5_7_7 : _GEN_561; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11367 = 3'h6 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11369 = 3'h6 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_563 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_6_0_0 : _GEN_562; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_564 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_6_0_1 : _GEN_563; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_565 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_6_0_2 : _GEN_564; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_566 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_6_0_3 : _GEN_565; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_567 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_6_0_4 : _GEN_566; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_568 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_6_0_5 : _GEN_567; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_569 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_6_0_6 : _GEN_568; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_570 = 3'h6 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_6_0_7 : _GEN_569; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11401 = 3'h6 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_571 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_6_1_0 : _GEN_570; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_572 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_6_1_1 : _GEN_571; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_573 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_6_1_2 : _GEN_572; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_574 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_6_1_3 : _GEN_573; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_575 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_6_1_4 : _GEN_574; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_576 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_6_1_5 : _GEN_575; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_577 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_6_1_6 : _GEN_576; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_578 = 3'h6 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_6_1_7 : _GEN_577; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11433 = 3'h6 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_579 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_6_2_0 : _GEN_578; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_580 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_6_2_1 : _GEN_579; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_581 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_6_2_2 : _GEN_580; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_582 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_6_2_3 : _GEN_581; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_583 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_6_2_4 : _GEN_582; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_584 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_6_2_5 : _GEN_583; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_585 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_6_2_6 : _GEN_584; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_586 = 3'h6 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_6_2_7 : _GEN_585; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11465 = 3'h6 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_587 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_6_3_0 : _GEN_586; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_588 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_6_3_1 : _GEN_587; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_589 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_6_3_2 : _GEN_588; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_590 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_6_3_3 : _GEN_589; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_591 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_6_3_4 : _GEN_590; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_592 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_6_3_5 : _GEN_591; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_593 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_6_3_6 : _GEN_592; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_594 = 3'h6 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_6_3_7 : _GEN_593; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11497 = 3'h6 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_595 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_6_4_0 : _GEN_594; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_596 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_6_4_1 : _GEN_595; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_597 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_6_4_2 : _GEN_596; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_598 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_6_4_3 : _GEN_597; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_599 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_6_4_4 : _GEN_598; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_600 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_6_4_5 : _GEN_599; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_601 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_6_4_6 : _GEN_600; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_602 = 3'h6 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_6_4_7 : _GEN_601; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11529 = 3'h6 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_603 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_6_5_0 : _GEN_602; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_604 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_6_5_1 : _GEN_603; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_605 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_6_5_2 : _GEN_604; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_606 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_6_5_3 : _GEN_605; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_607 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_6_5_4 : _GEN_606; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_608 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_6_5_5 : _GEN_607; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_609 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_6_5_6 : _GEN_608; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_610 = 3'h6 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_6_5_7 : _GEN_609; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11561 = 3'h6 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_611 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_6_6_0 : _GEN_610; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_612 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_6_6_1 : _GEN_611; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_613 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_6_6_2 : _GEN_612; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_614 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_6_6_3 : _GEN_613; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_615 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_6_6_4 : _GEN_614; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_616 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_6_6_5 : _GEN_615; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_617 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_6_6_6 : _GEN_616; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_618 = 3'h6 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_6_6_7 : _GEN_617; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11593 = 3'h6 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_619 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_6_7_0 : _GEN_618; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_620 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_6_7_1 : _GEN_619; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_621 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_6_7_2 : _GEN_620; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_622 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_6_7_3 : _GEN_621; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_623 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_6_7_4 : _GEN_622; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_624 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_6_7_5 : _GEN_623; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_625 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_6_7_6 : _GEN_624; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_626 = 3'h6 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_6_7_7 : _GEN_625; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11623 = 3'h7 == set_addr; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11625 = 3'h7 == set_addr & 3'h0 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_627 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h0 == line_addr ? CacheMem_7_0_0 : _GEN_626; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_628 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h1 == line_addr ? CacheMem_7_0_1 : _GEN_627; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_629 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h2 == line_addr ? CacheMem_7_0_2 : _GEN_628; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_630 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h3 == line_addr ? CacheMem_7_0_3 : _GEN_629; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_631 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h4 == line_addr ? CacheMem_7_0_4 : _GEN_630; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_632 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h5 == line_addr ? CacheMem_7_0_5 : _GEN_631; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_633 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h6 == line_addr ? CacheMem_7_0_6 : _GEN_632; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_634 = 3'h7 == set_addr & 3'h0 == way_hit & 3'h7 == line_addr ? CacheMem_7_0_7 : _GEN_633; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11657 = 3'h7 == set_addr & 3'h1 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_635 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h0 == line_addr ? CacheMem_7_1_0 : _GEN_634; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_636 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h1 == line_addr ? CacheMem_7_1_1 : _GEN_635; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_637 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h2 == line_addr ? CacheMem_7_1_2 : _GEN_636; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_638 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h3 == line_addr ? CacheMem_7_1_3 : _GEN_637; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_639 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h4 == line_addr ? CacheMem_7_1_4 : _GEN_638; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_640 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h5 == line_addr ? CacheMem_7_1_5 : _GEN_639; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_641 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h6 == line_addr ? CacheMem_7_1_6 : _GEN_640; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_642 = 3'h7 == set_addr & 3'h1 == way_hit & 3'h7 == line_addr ? CacheMem_7_1_7 : _GEN_641; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11689 = 3'h7 == set_addr & 3'h2 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_643 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h0 == line_addr ? CacheMem_7_2_0 : _GEN_642; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_644 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h1 == line_addr ? CacheMem_7_2_1 : _GEN_643; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_645 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h2 == line_addr ? CacheMem_7_2_2 : _GEN_644; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_646 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h3 == line_addr ? CacheMem_7_2_3 : _GEN_645; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_647 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h4 == line_addr ? CacheMem_7_2_4 : _GEN_646; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_648 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h5 == line_addr ? CacheMem_7_2_5 : _GEN_647; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_649 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h6 == line_addr ? CacheMem_7_2_6 : _GEN_648; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_650 = 3'h7 == set_addr & 3'h2 == way_hit & 3'h7 == line_addr ? CacheMem_7_2_7 : _GEN_649; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11721 = 3'h7 == set_addr & 3'h3 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_651 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h0 == line_addr ? CacheMem_7_3_0 : _GEN_650; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_652 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h1 == line_addr ? CacheMem_7_3_1 : _GEN_651; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_653 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h2 == line_addr ? CacheMem_7_3_2 : _GEN_652; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_654 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h3 == line_addr ? CacheMem_7_3_3 : _GEN_653; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_655 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h4 == line_addr ? CacheMem_7_3_4 : _GEN_654; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_656 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h5 == line_addr ? CacheMem_7_3_5 : _GEN_655; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_657 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h6 == line_addr ? CacheMem_7_3_6 : _GEN_656; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_658 = 3'h7 == set_addr & 3'h3 == way_hit & 3'h7 == line_addr ? CacheMem_7_3_7 : _GEN_657; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11753 = 3'h7 == set_addr & 3'h4 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_659 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h0 == line_addr ? CacheMem_7_4_0 : _GEN_658; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_660 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h1 == line_addr ? CacheMem_7_4_1 : _GEN_659; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_661 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h2 == line_addr ? CacheMem_7_4_2 : _GEN_660; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_662 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h3 == line_addr ? CacheMem_7_4_3 : _GEN_661; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_663 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h4 == line_addr ? CacheMem_7_4_4 : _GEN_662; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_664 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h5 == line_addr ? CacheMem_7_4_5 : _GEN_663; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_665 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h6 == line_addr ? CacheMem_7_4_6 : _GEN_664; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_666 = 3'h7 == set_addr & 3'h4 == way_hit & 3'h7 == line_addr ? CacheMem_7_4_7 : _GEN_665; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11785 = 3'h7 == set_addr & 3'h5 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_667 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h0 == line_addr ? CacheMem_7_5_0 : _GEN_666; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_668 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h1 == line_addr ? CacheMem_7_5_1 : _GEN_667; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_669 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h2 == line_addr ? CacheMem_7_5_2 : _GEN_668; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_670 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h3 == line_addr ? CacheMem_7_5_3 : _GEN_669; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_671 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h4 == line_addr ? CacheMem_7_5_4 : _GEN_670; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_672 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h5 == line_addr ? CacheMem_7_5_5 : _GEN_671; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_673 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h6 == line_addr ? CacheMem_7_5_6 : _GEN_672; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_674 = 3'h7 == set_addr & 3'h5 == way_hit & 3'h7 == line_addr ? CacheMem_7_5_7 : _GEN_673; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11817 = 3'h7 == set_addr & 3'h6 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_675 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h0 == line_addr ? CacheMem_7_6_0 : _GEN_674; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_676 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h1 == line_addr ? CacheMem_7_6_1 : _GEN_675; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_677 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h2 == line_addr ? CacheMem_7_6_2 : _GEN_676; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_678 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h3 == line_addr ? CacheMem_7_6_3 : _GEN_677; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_679 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h4 == line_addr ? CacheMem_7_6_4 : _GEN_678; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_680 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h5 == line_addr ? CacheMem_7_6_5 : _GEN_679; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_681 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h6 == line_addr ? CacheMem_7_6_6 : _GEN_680; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_682 = 3'h7 == set_addr & 3'h6 == way_hit & 3'h7 == line_addr ? CacheMem_7_6_7 : _GEN_681; // @[Cache.scala 131:{15,15}]
  wire  _GEN_11849 = 3'h7 == set_addr & 3'h7 == way_hit; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_683 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h0 == line_addr ? CacheMem_7_7_0 : _GEN_682; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_684 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h1 == line_addr ? CacheMem_7_7_1 : _GEN_683; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_685 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h2 == line_addr ? CacheMem_7_7_2 : _GEN_684; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_686 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h3 == line_addr ? CacheMem_7_7_3 : _GEN_685; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_687 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h4 == line_addr ? CacheMem_7_7_4 : _GEN_686; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_688 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h5 == line_addr ? CacheMem_7_7_5 : _GEN_687; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_689 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h6 == line_addr ? CacheMem_7_7_6 : _GEN_688; // @[Cache.scala 131:{15,15}]
  wire [31:0] _GEN_690 = 3'h7 == set_addr & 3'h7 == way_hit & 3'h7 == line_addr ? CacheMem_7_7_7 : _GEN_689; // @[Cache.scala 131:{15,15}]
  wire [31:0] _CacheMem_T_1 = {24'h0,io_writedata[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_691 = _GEN_9837 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_692 = _GEN_9837 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_693 = _GEN_9837 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_694 = _GEN_9837 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_695 = _GEN_9837 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_696 = _GEN_9837 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_697 = _GEN_9837 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_698 = _GEN_9837 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_699 = _GEN_9865 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_700 = _GEN_9865 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_701 = _GEN_9865 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_702 = _GEN_9865 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_703 = _GEN_9865 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_704 = _GEN_9865 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_705 = _GEN_9865 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_706 = _GEN_9865 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_707 = _GEN_9897 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_708 = _GEN_9897 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_709 = _GEN_9897 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_710 = _GEN_9897 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_711 = _GEN_9897 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_712 = _GEN_9897 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_713 = _GEN_9897 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_714 = _GEN_9897 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_715 = _GEN_9929 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_716 = _GEN_9929 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_717 = _GEN_9929 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_718 = _GEN_9929 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_719 = _GEN_9929 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_720 = _GEN_9929 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_721 = _GEN_9929 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_722 = _GEN_9929 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_723 = _GEN_9961 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_724 = _GEN_9961 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_725 = _GEN_9961 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_726 = _GEN_9961 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_727 = _GEN_9961 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_728 = _GEN_9961 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_729 = _GEN_9961 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_730 = _GEN_9961 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_731 = _GEN_9993 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_732 = _GEN_9993 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_733 = _GEN_9993 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_734 = _GEN_9993 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_735 = _GEN_9993 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_736 = _GEN_9993 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_737 = _GEN_9993 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_738 = _GEN_9993 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_739 = _GEN_10025 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_740 = _GEN_10025 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_741 = _GEN_10025 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_742 = _GEN_10025 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_743 = _GEN_10025 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_744 = _GEN_10025 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_745 = _GEN_10025 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_746 = _GEN_10025 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_747 = _GEN_10057 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_0_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_748 = _GEN_10057 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_0_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_749 = _GEN_10057 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_0_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_750 = _GEN_10057 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_0_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_751 = _GEN_10057 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_0_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_752 = _GEN_10057 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_0_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_753 = _GEN_10057 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_0_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_754 = _GEN_10057 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_0_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_755 = _GEN_10089 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_756 = _GEN_10089 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_757 = _GEN_10089 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_758 = _GEN_10089 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_759 = _GEN_10089 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_760 = _GEN_10089 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_761 = _GEN_10089 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_762 = _GEN_10089 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_763 = _GEN_10121 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_764 = _GEN_10121 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_765 = _GEN_10121 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_766 = _GEN_10121 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_767 = _GEN_10121 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_768 = _GEN_10121 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_769 = _GEN_10121 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_770 = _GEN_10121 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_771 = _GEN_10153 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_772 = _GEN_10153 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_773 = _GEN_10153 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_774 = _GEN_10153 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_775 = _GEN_10153 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_776 = _GEN_10153 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_777 = _GEN_10153 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_778 = _GEN_10153 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_779 = _GEN_10185 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_780 = _GEN_10185 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_781 = _GEN_10185 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_782 = _GEN_10185 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_783 = _GEN_10185 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_784 = _GEN_10185 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_785 = _GEN_10185 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_786 = _GEN_10185 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_787 = _GEN_10217 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_788 = _GEN_10217 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_789 = _GEN_10217 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_790 = _GEN_10217 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_791 = _GEN_10217 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_792 = _GEN_10217 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_793 = _GEN_10217 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_794 = _GEN_10217 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_795 = _GEN_10249 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_796 = _GEN_10249 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_797 = _GEN_10249 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_798 = _GEN_10249 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_799 = _GEN_10249 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_800 = _GEN_10249 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_801 = _GEN_10249 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_802 = _GEN_10249 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_803 = _GEN_10281 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_804 = _GEN_10281 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_805 = _GEN_10281 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_806 = _GEN_10281 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_807 = _GEN_10281 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_808 = _GEN_10281 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_809 = _GEN_10281 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_810 = _GEN_10281 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_811 = _GEN_10313 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_1_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_812 = _GEN_10313 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_1_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_813 = _GEN_10313 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_1_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_814 = _GEN_10313 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_1_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_815 = _GEN_10313 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_1_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_816 = _GEN_10313 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_1_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_817 = _GEN_10313 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_1_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_818 = _GEN_10313 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_1_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_819 = _GEN_10345 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_820 = _GEN_10345 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_821 = _GEN_10345 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_822 = _GEN_10345 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_823 = _GEN_10345 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_824 = _GEN_10345 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_825 = _GEN_10345 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_826 = _GEN_10345 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_827 = _GEN_10377 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_828 = _GEN_10377 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_829 = _GEN_10377 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_830 = _GEN_10377 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_831 = _GEN_10377 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_832 = _GEN_10377 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_833 = _GEN_10377 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_834 = _GEN_10377 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_835 = _GEN_10409 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_836 = _GEN_10409 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_837 = _GEN_10409 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_838 = _GEN_10409 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_839 = _GEN_10409 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_840 = _GEN_10409 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_841 = _GEN_10409 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_842 = _GEN_10409 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_843 = _GEN_10441 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_844 = _GEN_10441 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_845 = _GEN_10441 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_846 = _GEN_10441 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_847 = _GEN_10441 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_848 = _GEN_10441 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_849 = _GEN_10441 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_850 = _GEN_10441 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_851 = _GEN_10473 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_852 = _GEN_10473 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_853 = _GEN_10473 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_854 = _GEN_10473 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_855 = _GEN_10473 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_856 = _GEN_10473 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_857 = _GEN_10473 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_858 = _GEN_10473 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_859 = _GEN_10505 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_860 = _GEN_10505 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_861 = _GEN_10505 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_862 = _GEN_10505 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_863 = _GEN_10505 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_864 = _GEN_10505 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_865 = _GEN_10505 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_866 = _GEN_10505 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_867 = _GEN_10537 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_868 = _GEN_10537 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_869 = _GEN_10537 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_870 = _GEN_10537 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_871 = _GEN_10537 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_872 = _GEN_10537 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_873 = _GEN_10537 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_874 = _GEN_10537 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_875 = _GEN_10569 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_2_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_876 = _GEN_10569 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_2_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_877 = _GEN_10569 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_2_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_878 = _GEN_10569 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_2_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_879 = _GEN_10569 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_2_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_880 = _GEN_10569 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_2_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_881 = _GEN_10569 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_2_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_882 = _GEN_10569 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_2_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_883 = _GEN_10601 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_884 = _GEN_10601 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_885 = _GEN_10601 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_886 = _GEN_10601 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_887 = _GEN_10601 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_888 = _GEN_10601 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_889 = _GEN_10601 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_890 = _GEN_10601 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_891 = _GEN_10633 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_892 = _GEN_10633 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_893 = _GEN_10633 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_894 = _GEN_10633 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_895 = _GEN_10633 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_896 = _GEN_10633 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_897 = _GEN_10633 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_898 = _GEN_10633 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_899 = _GEN_10665 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_900 = _GEN_10665 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_901 = _GEN_10665 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_902 = _GEN_10665 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_903 = _GEN_10665 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_904 = _GEN_10665 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_905 = _GEN_10665 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_906 = _GEN_10665 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_907 = _GEN_10697 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_908 = _GEN_10697 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_909 = _GEN_10697 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_910 = _GEN_10697 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_911 = _GEN_10697 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_912 = _GEN_10697 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_913 = _GEN_10697 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_914 = _GEN_10697 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_915 = _GEN_10729 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_916 = _GEN_10729 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_917 = _GEN_10729 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_918 = _GEN_10729 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_919 = _GEN_10729 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_920 = _GEN_10729 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_921 = _GEN_10729 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_922 = _GEN_10729 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_923 = _GEN_10761 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_924 = _GEN_10761 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_925 = _GEN_10761 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_926 = _GEN_10761 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_927 = _GEN_10761 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_928 = _GEN_10761 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_929 = _GEN_10761 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_930 = _GEN_10761 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_931 = _GEN_10793 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_932 = _GEN_10793 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_933 = _GEN_10793 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_934 = _GEN_10793 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_935 = _GEN_10793 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_936 = _GEN_10793 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_937 = _GEN_10793 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_938 = _GEN_10793 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_939 = _GEN_10825 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_3_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_940 = _GEN_10825 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_3_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_941 = _GEN_10825 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_3_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_942 = _GEN_10825 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_3_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_943 = _GEN_10825 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_3_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_944 = _GEN_10825 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_3_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_945 = _GEN_10825 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_3_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_946 = _GEN_10825 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_3_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_947 = _GEN_10857 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_948 = _GEN_10857 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_949 = _GEN_10857 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_950 = _GEN_10857 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_951 = _GEN_10857 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_952 = _GEN_10857 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_953 = _GEN_10857 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_954 = _GEN_10857 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_955 = _GEN_10889 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_956 = _GEN_10889 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_957 = _GEN_10889 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_958 = _GEN_10889 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_959 = _GEN_10889 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_960 = _GEN_10889 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_961 = _GEN_10889 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_962 = _GEN_10889 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_963 = _GEN_10921 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_964 = _GEN_10921 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_965 = _GEN_10921 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_966 = _GEN_10921 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_967 = _GEN_10921 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_968 = _GEN_10921 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_969 = _GEN_10921 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_970 = _GEN_10921 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_971 = _GEN_10953 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_972 = _GEN_10953 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_973 = _GEN_10953 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_974 = _GEN_10953 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_975 = _GEN_10953 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_976 = _GEN_10953 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_977 = _GEN_10953 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_978 = _GEN_10953 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_979 = _GEN_10985 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_980 = _GEN_10985 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_981 = _GEN_10985 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_982 = _GEN_10985 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_983 = _GEN_10985 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_984 = _GEN_10985 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_985 = _GEN_10985 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_986 = _GEN_10985 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_987 = _GEN_11017 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_988 = _GEN_11017 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_989 = _GEN_11017 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_990 = _GEN_11017 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_991 = _GEN_11017 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_992 = _GEN_11017 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_993 = _GEN_11017 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_994 = _GEN_11017 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_995 = _GEN_11049 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_996 = _GEN_11049 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_997 = _GEN_11049 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_998 = _GEN_11049 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_999 = _GEN_11049 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1000 = _GEN_11049 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1001 = _GEN_11049 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1002 = _GEN_11049 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1003 = _GEN_11081 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_4_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1004 = _GEN_11081 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_4_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1005 = _GEN_11081 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_4_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1006 = _GEN_11081 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_4_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1007 = _GEN_11081 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_4_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1008 = _GEN_11081 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_4_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1009 = _GEN_11081 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_4_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1010 = _GEN_11081 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_4_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1011 = _GEN_11113 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1012 = _GEN_11113 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1013 = _GEN_11113 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1014 = _GEN_11113 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1015 = _GEN_11113 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1016 = _GEN_11113 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1017 = _GEN_11113 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1018 = _GEN_11113 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1019 = _GEN_11145 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1020 = _GEN_11145 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1021 = _GEN_11145 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1022 = _GEN_11145 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1023 = _GEN_11145 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1024 = _GEN_11145 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1025 = _GEN_11145 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1026 = _GEN_11145 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1027 = _GEN_11177 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1028 = _GEN_11177 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1029 = _GEN_11177 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1030 = _GEN_11177 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1031 = _GEN_11177 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1032 = _GEN_11177 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1033 = _GEN_11177 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1034 = _GEN_11177 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1035 = _GEN_11209 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1036 = _GEN_11209 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1037 = _GEN_11209 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1038 = _GEN_11209 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1039 = _GEN_11209 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1040 = _GEN_11209 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1041 = _GEN_11209 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1042 = _GEN_11209 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1043 = _GEN_11241 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1044 = _GEN_11241 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1045 = _GEN_11241 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1046 = _GEN_11241 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1047 = _GEN_11241 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1048 = _GEN_11241 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1049 = _GEN_11241 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1050 = _GEN_11241 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1051 = _GEN_11273 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1052 = _GEN_11273 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1053 = _GEN_11273 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1054 = _GEN_11273 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1055 = _GEN_11273 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1056 = _GEN_11273 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1057 = _GEN_11273 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1058 = _GEN_11273 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1059 = _GEN_11305 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1060 = _GEN_11305 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1061 = _GEN_11305 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1062 = _GEN_11305 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1063 = _GEN_11305 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1064 = _GEN_11305 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1065 = _GEN_11305 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1066 = _GEN_11305 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1067 = _GEN_11337 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_5_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1068 = _GEN_11337 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_5_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1069 = _GEN_11337 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_5_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1070 = _GEN_11337 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_5_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1071 = _GEN_11337 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_5_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1072 = _GEN_11337 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_5_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1073 = _GEN_11337 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_5_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1074 = _GEN_11337 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_5_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1075 = _GEN_11369 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1076 = _GEN_11369 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1077 = _GEN_11369 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1078 = _GEN_11369 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1079 = _GEN_11369 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1080 = _GEN_11369 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1081 = _GEN_11369 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1082 = _GEN_11369 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1083 = _GEN_11401 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1084 = _GEN_11401 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1085 = _GEN_11401 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1086 = _GEN_11401 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1087 = _GEN_11401 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1088 = _GEN_11401 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1089 = _GEN_11401 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1090 = _GEN_11401 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1091 = _GEN_11433 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1092 = _GEN_11433 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1093 = _GEN_11433 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1094 = _GEN_11433 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1095 = _GEN_11433 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1096 = _GEN_11433 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1097 = _GEN_11433 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1098 = _GEN_11433 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1099 = _GEN_11465 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1100 = _GEN_11465 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1101 = _GEN_11465 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1102 = _GEN_11465 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1103 = _GEN_11465 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1104 = _GEN_11465 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1105 = _GEN_11465 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1106 = _GEN_11465 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1107 = _GEN_11497 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1108 = _GEN_11497 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1109 = _GEN_11497 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1110 = _GEN_11497 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1111 = _GEN_11497 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1112 = _GEN_11497 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1113 = _GEN_11497 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1114 = _GEN_11497 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1115 = _GEN_11529 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1116 = _GEN_11529 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1117 = _GEN_11529 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1118 = _GEN_11529 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1119 = _GEN_11529 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1120 = _GEN_11529 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1121 = _GEN_11529 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1122 = _GEN_11529 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1123 = _GEN_11561 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1124 = _GEN_11561 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1125 = _GEN_11561 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1126 = _GEN_11561 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1127 = _GEN_11561 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1128 = _GEN_11561 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1129 = _GEN_11561 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1130 = _GEN_11561 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1131 = _GEN_11593 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_6_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1132 = _GEN_11593 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_6_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1133 = _GEN_11593 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_6_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1134 = _GEN_11593 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_6_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1135 = _GEN_11593 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_6_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1136 = _GEN_11593 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_6_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1137 = _GEN_11593 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_6_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1138 = _GEN_11593 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_6_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1139 = _GEN_11625 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_0_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1140 = _GEN_11625 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_0_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1141 = _GEN_11625 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_0_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1142 = _GEN_11625 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_0_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1143 = _GEN_11625 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_0_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1144 = _GEN_11625 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_0_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1145 = _GEN_11625 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_0_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1146 = _GEN_11625 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_0_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1147 = _GEN_11657 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_1_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1148 = _GEN_11657 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_1_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1149 = _GEN_11657 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_1_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1150 = _GEN_11657 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_1_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1151 = _GEN_11657 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_1_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1152 = _GEN_11657 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_1_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1153 = _GEN_11657 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_1_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1154 = _GEN_11657 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_1_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1155 = _GEN_11689 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_2_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1156 = _GEN_11689 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_2_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1157 = _GEN_11689 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_2_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1158 = _GEN_11689 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_2_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1159 = _GEN_11689 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_2_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1160 = _GEN_11689 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_2_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1161 = _GEN_11689 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_2_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1162 = _GEN_11689 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_2_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1163 = _GEN_11721 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_3_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1164 = _GEN_11721 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_3_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1165 = _GEN_11721 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_3_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1166 = _GEN_11721 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_3_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1167 = _GEN_11721 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_3_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1168 = _GEN_11721 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_3_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1169 = _GEN_11721 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_3_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1170 = _GEN_11721 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_3_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1171 = _GEN_11753 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_4_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1172 = _GEN_11753 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_4_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1173 = _GEN_11753 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_4_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1174 = _GEN_11753 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_4_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1175 = _GEN_11753 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_4_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1176 = _GEN_11753 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_4_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1177 = _GEN_11753 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_4_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1178 = _GEN_11753 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_4_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1179 = _GEN_11785 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_5_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1180 = _GEN_11785 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_5_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1181 = _GEN_11785 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_5_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1182 = _GEN_11785 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_5_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1183 = _GEN_11785 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_5_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1184 = _GEN_11785 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_5_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1185 = _GEN_11785 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_5_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1186 = _GEN_11785 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_5_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1187 = _GEN_11817 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_6_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1188 = _GEN_11817 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_6_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1189 = _GEN_11817 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_6_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1190 = _GEN_11817 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_6_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1191 = _GEN_11817 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_6_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1192 = _GEN_11817 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_6_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1193 = _GEN_11817 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_6_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1194 = _GEN_11817 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_6_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1195 = _GEN_11849 & _GEN_9866 ? _CacheMem_T_1 : CacheMem_7_7_0; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1196 = _GEN_11849 & _GEN_9838 ? _CacheMem_T_1 : CacheMem_7_7_1; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1197 = _GEN_11849 & _GEN_9842 ? _CacheMem_T_1 : CacheMem_7_7_2; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1198 = _GEN_11849 & _GEN_9846 ? _CacheMem_T_1 : CacheMem_7_7_3; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1199 = _GEN_11849 & _GEN_9850 ? _CacheMem_T_1 : CacheMem_7_7_4; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1200 = _GEN_11849 & _GEN_9854 ? _CacheMem_T_1 : CacheMem_7_7_5; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1201 = _GEN_11849 & _GEN_9858 ? _CacheMem_T_1 : CacheMem_7_7_6; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _GEN_1202 = _GEN_11849 & _GEN_9862 ? _CacheMem_T_1 : CacheMem_7_7_7; // @[Cache.scala 135:{54,54} 53:25]
  wire [31:0] _CacheMem_T_3 = {16'h0,io_writedata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_1203 = _GEN_9837 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1204 = _GEN_9837 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1205 = _GEN_9837 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1206 = _GEN_9837 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1207 = _GEN_9837 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1208 = _GEN_9837 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1209 = _GEN_9837 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1210 = _GEN_9837 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1211 = _GEN_9865 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1212 = _GEN_9865 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1213 = _GEN_9865 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1214 = _GEN_9865 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1215 = _GEN_9865 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1216 = _GEN_9865 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1217 = _GEN_9865 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1218 = _GEN_9865 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1219 = _GEN_9897 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1220 = _GEN_9897 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1221 = _GEN_9897 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1222 = _GEN_9897 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1223 = _GEN_9897 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1224 = _GEN_9897 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1225 = _GEN_9897 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1226 = _GEN_9897 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1227 = _GEN_9929 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1228 = _GEN_9929 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1229 = _GEN_9929 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1230 = _GEN_9929 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1231 = _GEN_9929 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1232 = _GEN_9929 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1233 = _GEN_9929 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1234 = _GEN_9929 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1235 = _GEN_9961 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1236 = _GEN_9961 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1237 = _GEN_9961 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1238 = _GEN_9961 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1239 = _GEN_9961 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1240 = _GEN_9961 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1241 = _GEN_9961 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1242 = _GEN_9961 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1243 = _GEN_9993 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1244 = _GEN_9993 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1245 = _GEN_9993 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1246 = _GEN_9993 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1247 = _GEN_9993 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1248 = _GEN_9993 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1249 = _GEN_9993 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1250 = _GEN_9993 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1251 = _GEN_10025 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1252 = _GEN_10025 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1253 = _GEN_10025 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1254 = _GEN_10025 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1255 = _GEN_10025 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1256 = _GEN_10025 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1257 = _GEN_10025 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1258 = _GEN_10025 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1259 = _GEN_10057 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_0_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1260 = _GEN_10057 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_0_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1261 = _GEN_10057 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_0_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1262 = _GEN_10057 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_0_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1263 = _GEN_10057 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_0_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1264 = _GEN_10057 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_0_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1265 = _GEN_10057 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_0_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1266 = _GEN_10057 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_0_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1267 = _GEN_10089 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1268 = _GEN_10089 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1269 = _GEN_10089 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1270 = _GEN_10089 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1271 = _GEN_10089 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1272 = _GEN_10089 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1273 = _GEN_10089 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1274 = _GEN_10089 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1275 = _GEN_10121 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1276 = _GEN_10121 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1277 = _GEN_10121 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1278 = _GEN_10121 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1279 = _GEN_10121 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1280 = _GEN_10121 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1281 = _GEN_10121 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1282 = _GEN_10121 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1283 = _GEN_10153 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1284 = _GEN_10153 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1285 = _GEN_10153 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1286 = _GEN_10153 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1287 = _GEN_10153 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1288 = _GEN_10153 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1289 = _GEN_10153 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1290 = _GEN_10153 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1291 = _GEN_10185 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1292 = _GEN_10185 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1293 = _GEN_10185 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1294 = _GEN_10185 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1295 = _GEN_10185 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1296 = _GEN_10185 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1297 = _GEN_10185 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1298 = _GEN_10185 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1299 = _GEN_10217 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1300 = _GEN_10217 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1301 = _GEN_10217 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1302 = _GEN_10217 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1303 = _GEN_10217 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1304 = _GEN_10217 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1305 = _GEN_10217 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1306 = _GEN_10217 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1307 = _GEN_10249 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1308 = _GEN_10249 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1309 = _GEN_10249 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1310 = _GEN_10249 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1311 = _GEN_10249 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1312 = _GEN_10249 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1313 = _GEN_10249 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1314 = _GEN_10249 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1315 = _GEN_10281 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1316 = _GEN_10281 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1317 = _GEN_10281 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1318 = _GEN_10281 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1319 = _GEN_10281 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1320 = _GEN_10281 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1321 = _GEN_10281 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1322 = _GEN_10281 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1323 = _GEN_10313 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_1_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1324 = _GEN_10313 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_1_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1325 = _GEN_10313 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_1_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1326 = _GEN_10313 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_1_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1327 = _GEN_10313 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_1_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1328 = _GEN_10313 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_1_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1329 = _GEN_10313 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_1_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1330 = _GEN_10313 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_1_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1331 = _GEN_10345 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1332 = _GEN_10345 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1333 = _GEN_10345 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1334 = _GEN_10345 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1335 = _GEN_10345 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1336 = _GEN_10345 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1337 = _GEN_10345 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1338 = _GEN_10345 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1339 = _GEN_10377 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1340 = _GEN_10377 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1341 = _GEN_10377 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1342 = _GEN_10377 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1343 = _GEN_10377 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1344 = _GEN_10377 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1345 = _GEN_10377 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1346 = _GEN_10377 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1347 = _GEN_10409 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1348 = _GEN_10409 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1349 = _GEN_10409 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1350 = _GEN_10409 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1351 = _GEN_10409 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1352 = _GEN_10409 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1353 = _GEN_10409 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1354 = _GEN_10409 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1355 = _GEN_10441 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1356 = _GEN_10441 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1357 = _GEN_10441 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1358 = _GEN_10441 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1359 = _GEN_10441 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1360 = _GEN_10441 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1361 = _GEN_10441 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1362 = _GEN_10441 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1363 = _GEN_10473 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1364 = _GEN_10473 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1365 = _GEN_10473 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1366 = _GEN_10473 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1367 = _GEN_10473 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1368 = _GEN_10473 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1369 = _GEN_10473 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1370 = _GEN_10473 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1371 = _GEN_10505 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1372 = _GEN_10505 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1373 = _GEN_10505 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1374 = _GEN_10505 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1375 = _GEN_10505 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1376 = _GEN_10505 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1377 = _GEN_10505 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1378 = _GEN_10505 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1379 = _GEN_10537 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1380 = _GEN_10537 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1381 = _GEN_10537 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1382 = _GEN_10537 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1383 = _GEN_10537 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1384 = _GEN_10537 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1385 = _GEN_10537 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1386 = _GEN_10537 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1387 = _GEN_10569 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_2_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1388 = _GEN_10569 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_2_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1389 = _GEN_10569 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_2_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1390 = _GEN_10569 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_2_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1391 = _GEN_10569 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_2_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1392 = _GEN_10569 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_2_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1393 = _GEN_10569 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_2_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1394 = _GEN_10569 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_2_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1395 = _GEN_10601 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1396 = _GEN_10601 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1397 = _GEN_10601 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1398 = _GEN_10601 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1399 = _GEN_10601 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1400 = _GEN_10601 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1401 = _GEN_10601 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1402 = _GEN_10601 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1403 = _GEN_10633 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1404 = _GEN_10633 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1405 = _GEN_10633 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1406 = _GEN_10633 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1407 = _GEN_10633 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1408 = _GEN_10633 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1409 = _GEN_10633 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1410 = _GEN_10633 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1411 = _GEN_10665 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1412 = _GEN_10665 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1413 = _GEN_10665 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1414 = _GEN_10665 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1415 = _GEN_10665 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1416 = _GEN_10665 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1417 = _GEN_10665 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1418 = _GEN_10665 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1419 = _GEN_10697 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1420 = _GEN_10697 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1421 = _GEN_10697 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1422 = _GEN_10697 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1423 = _GEN_10697 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1424 = _GEN_10697 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1425 = _GEN_10697 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1426 = _GEN_10697 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1427 = _GEN_10729 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1428 = _GEN_10729 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1429 = _GEN_10729 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1430 = _GEN_10729 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1431 = _GEN_10729 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1432 = _GEN_10729 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1433 = _GEN_10729 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1434 = _GEN_10729 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1435 = _GEN_10761 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1436 = _GEN_10761 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1437 = _GEN_10761 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1438 = _GEN_10761 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1439 = _GEN_10761 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1440 = _GEN_10761 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1441 = _GEN_10761 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1442 = _GEN_10761 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1443 = _GEN_10793 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1444 = _GEN_10793 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1445 = _GEN_10793 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1446 = _GEN_10793 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1447 = _GEN_10793 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1448 = _GEN_10793 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1449 = _GEN_10793 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1450 = _GEN_10793 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1451 = _GEN_10825 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_3_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1452 = _GEN_10825 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_3_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1453 = _GEN_10825 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_3_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1454 = _GEN_10825 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_3_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1455 = _GEN_10825 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_3_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1456 = _GEN_10825 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_3_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1457 = _GEN_10825 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_3_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1458 = _GEN_10825 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_3_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1459 = _GEN_10857 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1460 = _GEN_10857 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1461 = _GEN_10857 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1462 = _GEN_10857 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1463 = _GEN_10857 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1464 = _GEN_10857 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1465 = _GEN_10857 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1466 = _GEN_10857 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1467 = _GEN_10889 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1468 = _GEN_10889 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1469 = _GEN_10889 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1470 = _GEN_10889 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1471 = _GEN_10889 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1472 = _GEN_10889 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1473 = _GEN_10889 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1474 = _GEN_10889 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1475 = _GEN_10921 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1476 = _GEN_10921 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1477 = _GEN_10921 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1478 = _GEN_10921 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1479 = _GEN_10921 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1480 = _GEN_10921 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1481 = _GEN_10921 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1482 = _GEN_10921 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1483 = _GEN_10953 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1484 = _GEN_10953 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1485 = _GEN_10953 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1486 = _GEN_10953 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1487 = _GEN_10953 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1488 = _GEN_10953 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1489 = _GEN_10953 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1490 = _GEN_10953 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1491 = _GEN_10985 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1492 = _GEN_10985 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1493 = _GEN_10985 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1494 = _GEN_10985 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1495 = _GEN_10985 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1496 = _GEN_10985 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1497 = _GEN_10985 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1498 = _GEN_10985 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1499 = _GEN_11017 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1500 = _GEN_11017 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1501 = _GEN_11017 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1502 = _GEN_11017 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1503 = _GEN_11017 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1504 = _GEN_11017 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1505 = _GEN_11017 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1506 = _GEN_11017 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1507 = _GEN_11049 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1508 = _GEN_11049 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1509 = _GEN_11049 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1510 = _GEN_11049 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1511 = _GEN_11049 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1512 = _GEN_11049 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1513 = _GEN_11049 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1514 = _GEN_11049 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1515 = _GEN_11081 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_4_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1516 = _GEN_11081 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_4_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1517 = _GEN_11081 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_4_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1518 = _GEN_11081 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_4_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1519 = _GEN_11081 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_4_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1520 = _GEN_11081 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_4_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1521 = _GEN_11081 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_4_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1522 = _GEN_11081 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_4_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1523 = _GEN_11113 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1524 = _GEN_11113 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1525 = _GEN_11113 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1526 = _GEN_11113 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1527 = _GEN_11113 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1528 = _GEN_11113 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1529 = _GEN_11113 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1530 = _GEN_11113 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1531 = _GEN_11145 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1532 = _GEN_11145 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1533 = _GEN_11145 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1534 = _GEN_11145 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1535 = _GEN_11145 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1536 = _GEN_11145 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1537 = _GEN_11145 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1538 = _GEN_11145 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1539 = _GEN_11177 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1540 = _GEN_11177 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1541 = _GEN_11177 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1542 = _GEN_11177 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1543 = _GEN_11177 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1544 = _GEN_11177 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1545 = _GEN_11177 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1546 = _GEN_11177 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1547 = _GEN_11209 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1548 = _GEN_11209 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1549 = _GEN_11209 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1550 = _GEN_11209 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1551 = _GEN_11209 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1552 = _GEN_11209 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1553 = _GEN_11209 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1554 = _GEN_11209 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1555 = _GEN_11241 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1556 = _GEN_11241 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1557 = _GEN_11241 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1558 = _GEN_11241 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1559 = _GEN_11241 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1560 = _GEN_11241 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1561 = _GEN_11241 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1562 = _GEN_11241 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1563 = _GEN_11273 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1564 = _GEN_11273 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1565 = _GEN_11273 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1566 = _GEN_11273 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1567 = _GEN_11273 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1568 = _GEN_11273 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1569 = _GEN_11273 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1570 = _GEN_11273 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1571 = _GEN_11305 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1572 = _GEN_11305 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1573 = _GEN_11305 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1574 = _GEN_11305 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1575 = _GEN_11305 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1576 = _GEN_11305 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1577 = _GEN_11305 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1578 = _GEN_11305 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1579 = _GEN_11337 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_5_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1580 = _GEN_11337 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_5_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1581 = _GEN_11337 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_5_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1582 = _GEN_11337 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_5_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1583 = _GEN_11337 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_5_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1584 = _GEN_11337 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_5_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1585 = _GEN_11337 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_5_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1586 = _GEN_11337 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_5_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1587 = _GEN_11369 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1588 = _GEN_11369 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1589 = _GEN_11369 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1590 = _GEN_11369 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1591 = _GEN_11369 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1592 = _GEN_11369 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1593 = _GEN_11369 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1594 = _GEN_11369 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1595 = _GEN_11401 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1596 = _GEN_11401 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1597 = _GEN_11401 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1598 = _GEN_11401 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1599 = _GEN_11401 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1600 = _GEN_11401 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1601 = _GEN_11401 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1602 = _GEN_11401 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1603 = _GEN_11433 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1604 = _GEN_11433 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1605 = _GEN_11433 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1606 = _GEN_11433 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1607 = _GEN_11433 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1608 = _GEN_11433 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1609 = _GEN_11433 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1610 = _GEN_11433 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1611 = _GEN_11465 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1612 = _GEN_11465 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1613 = _GEN_11465 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1614 = _GEN_11465 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1615 = _GEN_11465 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1616 = _GEN_11465 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1617 = _GEN_11465 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1618 = _GEN_11465 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1619 = _GEN_11497 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1620 = _GEN_11497 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1621 = _GEN_11497 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1622 = _GEN_11497 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1623 = _GEN_11497 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1624 = _GEN_11497 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1625 = _GEN_11497 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1626 = _GEN_11497 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1627 = _GEN_11529 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1628 = _GEN_11529 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1629 = _GEN_11529 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1630 = _GEN_11529 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1631 = _GEN_11529 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1632 = _GEN_11529 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1633 = _GEN_11529 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1634 = _GEN_11529 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1635 = _GEN_11561 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1636 = _GEN_11561 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1637 = _GEN_11561 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1638 = _GEN_11561 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1639 = _GEN_11561 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1640 = _GEN_11561 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1641 = _GEN_11561 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1642 = _GEN_11561 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1643 = _GEN_11593 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_6_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1644 = _GEN_11593 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_6_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1645 = _GEN_11593 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_6_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1646 = _GEN_11593 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_6_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1647 = _GEN_11593 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_6_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1648 = _GEN_11593 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_6_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1649 = _GEN_11593 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_6_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1650 = _GEN_11593 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_6_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1651 = _GEN_11625 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_0_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1652 = _GEN_11625 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_0_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1653 = _GEN_11625 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_0_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1654 = _GEN_11625 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_0_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1655 = _GEN_11625 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_0_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1656 = _GEN_11625 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_0_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1657 = _GEN_11625 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_0_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1658 = _GEN_11625 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_0_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1659 = _GEN_11657 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_1_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1660 = _GEN_11657 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_1_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1661 = _GEN_11657 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_1_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1662 = _GEN_11657 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_1_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1663 = _GEN_11657 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_1_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1664 = _GEN_11657 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_1_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1665 = _GEN_11657 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_1_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1666 = _GEN_11657 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_1_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1667 = _GEN_11689 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_2_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1668 = _GEN_11689 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_2_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1669 = _GEN_11689 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_2_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1670 = _GEN_11689 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_2_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1671 = _GEN_11689 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_2_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1672 = _GEN_11689 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_2_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1673 = _GEN_11689 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_2_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1674 = _GEN_11689 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_2_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1675 = _GEN_11721 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_3_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1676 = _GEN_11721 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_3_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1677 = _GEN_11721 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_3_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1678 = _GEN_11721 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_3_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1679 = _GEN_11721 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_3_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1680 = _GEN_11721 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_3_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1681 = _GEN_11721 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_3_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1682 = _GEN_11721 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_3_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1683 = _GEN_11753 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_4_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1684 = _GEN_11753 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_4_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1685 = _GEN_11753 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_4_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1686 = _GEN_11753 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_4_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1687 = _GEN_11753 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_4_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1688 = _GEN_11753 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_4_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1689 = _GEN_11753 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_4_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1690 = _GEN_11753 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_4_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1691 = _GEN_11785 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_5_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1692 = _GEN_11785 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_5_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1693 = _GEN_11785 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_5_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1694 = _GEN_11785 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_5_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1695 = _GEN_11785 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_5_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1696 = _GEN_11785 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_5_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1697 = _GEN_11785 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_5_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1698 = _GEN_11785 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_5_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1699 = _GEN_11817 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_6_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1700 = _GEN_11817 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_6_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1701 = _GEN_11817 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_6_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1702 = _GEN_11817 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_6_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1703 = _GEN_11817 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_6_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1704 = _GEN_11817 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_6_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1705 = _GEN_11817 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_6_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1706 = _GEN_11817 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_6_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1707 = _GEN_11849 & _GEN_9866 ? _CacheMem_T_3 : CacheMem_7_7_0; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1708 = _GEN_11849 & _GEN_9838 ? _CacheMem_T_3 : CacheMem_7_7_1; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1709 = _GEN_11849 & _GEN_9842 ? _CacheMem_T_3 : CacheMem_7_7_2; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1710 = _GEN_11849 & _GEN_9846 ? _CacheMem_T_3 : CacheMem_7_7_3; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1711 = _GEN_11849 & _GEN_9850 ? _CacheMem_T_3 : CacheMem_7_7_4; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1712 = _GEN_11849 & _GEN_9854 ? _CacheMem_T_3 : CacheMem_7_7_5; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1713 = _GEN_11849 & _GEN_9858 ? _CacheMem_T_3 : CacheMem_7_7_6; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1714 = _GEN_11849 & _GEN_9862 ? _CacheMem_T_3 : CacheMem_7_7_7; // @[Cache.scala 138:{54,54} 53:25]
  wire [31:0] _GEN_1715 = _GEN_9837 & _GEN_9866 ? io_writedata : CacheMem_0_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1716 = _GEN_9837 & _GEN_9838 ? io_writedata : CacheMem_0_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1717 = _GEN_9837 & _GEN_9842 ? io_writedata : CacheMem_0_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1718 = _GEN_9837 & _GEN_9846 ? io_writedata : CacheMem_0_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1719 = _GEN_9837 & _GEN_9850 ? io_writedata : CacheMem_0_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1720 = _GEN_9837 & _GEN_9854 ? io_writedata : CacheMem_0_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1721 = _GEN_9837 & _GEN_9858 ? io_writedata : CacheMem_0_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1722 = _GEN_9837 & _GEN_9862 ? io_writedata : CacheMem_0_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1723 = _GEN_9865 & _GEN_9866 ? io_writedata : CacheMem_0_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1724 = _GEN_9865 & _GEN_9838 ? io_writedata : CacheMem_0_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1725 = _GEN_9865 & _GEN_9842 ? io_writedata : CacheMem_0_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1726 = _GEN_9865 & _GEN_9846 ? io_writedata : CacheMem_0_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1727 = _GEN_9865 & _GEN_9850 ? io_writedata : CacheMem_0_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1728 = _GEN_9865 & _GEN_9854 ? io_writedata : CacheMem_0_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1729 = _GEN_9865 & _GEN_9858 ? io_writedata : CacheMem_0_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1730 = _GEN_9865 & _GEN_9862 ? io_writedata : CacheMem_0_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1731 = _GEN_9897 & _GEN_9866 ? io_writedata : CacheMem_0_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1732 = _GEN_9897 & _GEN_9838 ? io_writedata : CacheMem_0_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1733 = _GEN_9897 & _GEN_9842 ? io_writedata : CacheMem_0_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1734 = _GEN_9897 & _GEN_9846 ? io_writedata : CacheMem_0_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1735 = _GEN_9897 & _GEN_9850 ? io_writedata : CacheMem_0_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1736 = _GEN_9897 & _GEN_9854 ? io_writedata : CacheMem_0_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1737 = _GEN_9897 & _GEN_9858 ? io_writedata : CacheMem_0_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1738 = _GEN_9897 & _GEN_9862 ? io_writedata : CacheMem_0_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1739 = _GEN_9929 & _GEN_9866 ? io_writedata : CacheMem_0_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1740 = _GEN_9929 & _GEN_9838 ? io_writedata : CacheMem_0_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1741 = _GEN_9929 & _GEN_9842 ? io_writedata : CacheMem_0_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1742 = _GEN_9929 & _GEN_9846 ? io_writedata : CacheMem_0_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1743 = _GEN_9929 & _GEN_9850 ? io_writedata : CacheMem_0_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1744 = _GEN_9929 & _GEN_9854 ? io_writedata : CacheMem_0_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1745 = _GEN_9929 & _GEN_9858 ? io_writedata : CacheMem_0_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1746 = _GEN_9929 & _GEN_9862 ? io_writedata : CacheMem_0_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1747 = _GEN_9961 & _GEN_9866 ? io_writedata : CacheMem_0_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1748 = _GEN_9961 & _GEN_9838 ? io_writedata : CacheMem_0_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1749 = _GEN_9961 & _GEN_9842 ? io_writedata : CacheMem_0_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1750 = _GEN_9961 & _GEN_9846 ? io_writedata : CacheMem_0_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1751 = _GEN_9961 & _GEN_9850 ? io_writedata : CacheMem_0_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1752 = _GEN_9961 & _GEN_9854 ? io_writedata : CacheMem_0_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1753 = _GEN_9961 & _GEN_9858 ? io_writedata : CacheMem_0_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1754 = _GEN_9961 & _GEN_9862 ? io_writedata : CacheMem_0_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1755 = _GEN_9993 & _GEN_9866 ? io_writedata : CacheMem_0_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1756 = _GEN_9993 & _GEN_9838 ? io_writedata : CacheMem_0_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1757 = _GEN_9993 & _GEN_9842 ? io_writedata : CacheMem_0_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1758 = _GEN_9993 & _GEN_9846 ? io_writedata : CacheMem_0_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1759 = _GEN_9993 & _GEN_9850 ? io_writedata : CacheMem_0_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1760 = _GEN_9993 & _GEN_9854 ? io_writedata : CacheMem_0_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1761 = _GEN_9993 & _GEN_9858 ? io_writedata : CacheMem_0_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1762 = _GEN_9993 & _GEN_9862 ? io_writedata : CacheMem_0_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1763 = _GEN_10025 & _GEN_9866 ? io_writedata : CacheMem_0_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1764 = _GEN_10025 & _GEN_9838 ? io_writedata : CacheMem_0_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1765 = _GEN_10025 & _GEN_9842 ? io_writedata : CacheMem_0_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1766 = _GEN_10025 & _GEN_9846 ? io_writedata : CacheMem_0_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1767 = _GEN_10025 & _GEN_9850 ? io_writedata : CacheMem_0_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1768 = _GEN_10025 & _GEN_9854 ? io_writedata : CacheMem_0_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1769 = _GEN_10025 & _GEN_9858 ? io_writedata : CacheMem_0_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1770 = _GEN_10025 & _GEN_9862 ? io_writedata : CacheMem_0_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1771 = _GEN_10057 & _GEN_9866 ? io_writedata : CacheMem_0_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1772 = _GEN_10057 & _GEN_9838 ? io_writedata : CacheMem_0_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1773 = _GEN_10057 & _GEN_9842 ? io_writedata : CacheMem_0_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1774 = _GEN_10057 & _GEN_9846 ? io_writedata : CacheMem_0_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1775 = _GEN_10057 & _GEN_9850 ? io_writedata : CacheMem_0_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1776 = _GEN_10057 & _GEN_9854 ? io_writedata : CacheMem_0_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1777 = _GEN_10057 & _GEN_9858 ? io_writedata : CacheMem_0_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1778 = _GEN_10057 & _GEN_9862 ? io_writedata : CacheMem_0_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1779 = _GEN_10089 & _GEN_9866 ? io_writedata : CacheMem_1_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1780 = _GEN_10089 & _GEN_9838 ? io_writedata : CacheMem_1_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1781 = _GEN_10089 & _GEN_9842 ? io_writedata : CacheMem_1_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1782 = _GEN_10089 & _GEN_9846 ? io_writedata : CacheMem_1_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1783 = _GEN_10089 & _GEN_9850 ? io_writedata : CacheMem_1_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1784 = _GEN_10089 & _GEN_9854 ? io_writedata : CacheMem_1_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1785 = _GEN_10089 & _GEN_9858 ? io_writedata : CacheMem_1_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1786 = _GEN_10089 & _GEN_9862 ? io_writedata : CacheMem_1_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1787 = _GEN_10121 & _GEN_9866 ? io_writedata : CacheMem_1_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1788 = _GEN_10121 & _GEN_9838 ? io_writedata : CacheMem_1_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1789 = _GEN_10121 & _GEN_9842 ? io_writedata : CacheMem_1_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1790 = _GEN_10121 & _GEN_9846 ? io_writedata : CacheMem_1_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1791 = _GEN_10121 & _GEN_9850 ? io_writedata : CacheMem_1_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1792 = _GEN_10121 & _GEN_9854 ? io_writedata : CacheMem_1_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1793 = _GEN_10121 & _GEN_9858 ? io_writedata : CacheMem_1_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1794 = _GEN_10121 & _GEN_9862 ? io_writedata : CacheMem_1_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1795 = _GEN_10153 & _GEN_9866 ? io_writedata : CacheMem_1_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1796 = _GEN_10153 & _GEN_9838 ? io_writedata : CacheMem_1_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1797 = _GEN_10153 & _GEN_9842 ? io_writedata : CacheMem_1_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1798 = _GEN_10153 & _GEN_9846 ? io_writedata : CacheMem_1_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1799 = _GEN_10153 & _GEN_9850 ? io_writedata : CacheMem_1_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1800 = _GEN_10153 & _GEN_9854 ? io_writedata : CacheMem_1_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1801 = _GEN_10153 & _GEN_9858 ? io_writedata : CacheMem_1_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1802 = _GEN_10153 & _GEN_9862 ? io_writedata : CacheMem_1_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1803 = _GEN_10185 & _GEN_9866 ? io_writedata : CacheMem_1_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1804 = _GEN_10185 & _GEN_9838 ? io_writedata : CacheMem_1_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1805 = _GEN_10185 & _GEN_9842 ? io_writedata : CacheMem_1_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1806 = _GEN_10185 & _GEN_9846 ? io_writedata : CacheMem_1_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1807 = _GEN_10185 & _GEN_9850 ? io_writedata : CacheMem_1_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1808 = _GEN_10185 & _GEN_9854 ? io_writedata : CacheMem_1_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1809 = _GEN_10185 & _GEN_9858 ? io_writedata : CacheMem_1_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1810 = _GEN_10185 & _GEN_9862 ? io_writedata : CacheMem_1_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1811 = _GEN_10217 & _GEN_9866 ? io_writedata : CacheMem_1_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1812 = _GEN_10217 & _GEN_9838 ? io_writedata : CacheMem_1_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1813 = _GEN_10217 & _GEN_9842 ? io_writedata : CacheMem_1_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1814 = _GEN_10217 & _GEN_9846 ? io_writedata : CacheMem_1_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1815 = _GEN_10217 & _GEN_9850 ? io_writedata : CacheMem_1_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1816 = _GEN_10217 & _GEN_9854 ? io_writedata : CacheMem_1_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1817 = _GEN_10217 & _GEN_9858 ? io_writedata : CacheMem_1_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1818 = _GEN_10217 & _GEN_9862 ? io_writedata : CacheMem_1_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1819 = _GEN_10249 & _GEN_9866 ? io_writedata : CacheMem_1_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1820 = _GEN_10249 & _GEN_9838 ? io_writedata : CacheMem_1_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1821 = _GEN_10249 & _GEN_9842 ? io_writedata : CacheMem_1_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1822 = _GEN_10249 & _GEN_9846 ? io_writedata : CacheMem_1_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1823 = _GEN_10249 & _GEN_9850 ? io_writedata : CacheMem_1_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1824 = _GEN_10249 & _GEN_9854 ? io_writedata : CacheMem_1_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1825 = _GEN_10249 & _GEN_9858 ? io_writedata : CacheMem_1_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1826 = _GEN_10249 & _GEN_9862 ? io_writedata : CacheMem_1_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1827 = _GEN_10281 & _GEN_9866 ? io_writedata : CacheMem_1_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1828 = _GEN_10281 & _GEN_9838 ? io_writedata : CacheMem_1_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1829 = _GEN_10281 & _GEN_9842 ? io_writedata : CacheMem_1_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1830 = _GEN_10281 & _GEN_9846 ? io_writedata : CacheMem_1_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1831 = _GEN_10281 & _GEN_9850 ? io_writedata : CacheMem_1_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1832 = _GEN_10281 & _GEN_9854 ? io_writedata : CacheMem_1_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1833 = _GEN_10281 & _GEN_9858 ? io_writedata : CacheMem_1_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1834 = _GEN_10281 & _GEN_9862 ? io_writedata : CacheMem_1_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1835 = _GEN_10313 & _GEN_9866 ? io_writedata : CacheMem_1_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1836 = _GEN_10313 & _GEN_9838 ? io_writedata : CacheMem_1_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1837 = _GEN_10313 & _GEN_9842 ? io_writedata : CacheMem_1_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1838 = _GEN_10313 & _GEN_9846 ? io_writedata : CacheMem_1_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1839 = _GEN_10313 & _GEN_9850 ? io_writedata : CacheMem_1_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1840 = _GEN_10313 & _GEN_9854 ? io_writedata : CacheMem_1_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1841 = _GEN_10313 & _GEN_9858 ? io_writedata : CacheMem_1_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1842 = _GEN_10313 & _GEN_9862 ? io_writedata : CacheMem_1_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1843 = _GEN_10345 & _GEN_9866 ? io_writedata : CacheMem_2_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1844 = _GEN_10345 & _GEN_9838 ? io_writedata : CacheMem_2_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1845 = _GEN_10345 & _GEN_9842 ? io_writedata : CacheMem_2_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1846 = _GEN_10345 & _GEN_9846 ? io_writedata : CacheMem_2_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1847 = _GEN_10345 & _GEN_9850 ? io_writedata : CacheMem_2_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1848 = _GEN_10345 & _GEN_9854 ? io_writedata : CacheMem_2_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1849 = _GEN_10345 & _GEN_9858 ? io_writedata : CacheMem_2_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1850 = _GEN_10345 & _GEN_9862 ? io_writedata : CacheMem_2_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1851 = _GEN_10377 & _GEN_9866 ? io_writedata : CacheMem_2_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1852 = _GEN_10377 & _GEN_9838 ? io_writedata : CacheMem_2_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1853 = _GEN_10377 & _GEN_9842 ? io_writedata : CacheMem_2_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1854 = _GEN_10377 & _GEN_9846 ? io_writedata : CacheMem_2_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1855 = _GEN_10377 & _GEN_9850 ? io_writedata : CacheMem_2_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1856 = _GEN_10377 & _GEN_9854 ? io_writedata : CacheMem_2_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1857 = _GEN_10377 & _GEN_9858 ? io_writedata : CacheMem_2_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1858 = _GEN_10377 & _GEN_9862 ? io_writedata : CacheMem_2_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1859 = _GEN_10409 & _GEN_9866 ? io_writedata : CacheMem_2_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1860 = _GEN_10409 & _GEN_9838 ? io_writedata : CacheMem_2_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1861 = _GEN_10409 & _GEN_9842 ? io_writedata : CacheMem_2_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1862 = _GEN_10409 & _GEN_9846 ? io_writedata : CacheMem_2_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1863 = _GEN_10409 & _GEN_9850 ? io_writedata : CacheMem_2_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1864 = _GEN_10409 & _GEN_9854 ? io_writedata : CacheMem_2_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1865 = _GEN_10409 & _GEN_9858 ? io_writedata : CacheMem_2_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1866 = _GEN_10409 & _GEN_9862 ? io_writedata : CacheMem_2_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1867 = _GEN_10441 & _GEN_9866 ? io_writedata : CacheMem_2_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1868 = _GEN_10441 & _GEN_9838 ? io_writedata : CacheMem_2_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1869 = _GEN_10441 & _GEN_9842 ? io_writedata : CacheMem_2_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1870 = _GEN_10441 & _GEN_9846 ? io_writedata : CacheMem_2_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1871 = _GEN_10441 & _GEN_9850 ? io_writedata : CacheMem_2_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1872 = _GEN_10441 & _GEN_9854 ? io_writedata : CacheMem_2_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1873 = _GEN_10441 & _GEN_9858 ? io_writedata : CacheMem_2_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1874 = _GEN_10441 & _GEN_9862 ? io_writedata : CacheMem_2_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1875 = _GEN_10473 & _GEN_9866 ? io_writedata : CacheMem_2_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1876 = _GEN_10473 & _GEN_9838 ? io_writedata : CacheMem_2_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1877 = _GEN_10473 & _GEN_9842 ? io_writedata : CacheMem_2_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1878 = _GEN_10473 & _GEN_9846 ? io_writedata : CacheMem_2_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1879 = _GEN_10473 & _GEN_9850 ? io_writedata : CacheMem_2_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1880 = _GEN_10473 & _GEN_9854 ? io_writedata : CacheMem_2_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1881 = _GEN_10473 & _GEN_9858 ? io_writedata : CacheMem_2_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1882 = _GEN_10473 & _GEN_9862 ? io_writedata : CacheMem_2_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1883 = _GEN_10505 & _GEN_9866 ? io_writedata : CacheMem_2_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1884 = _GEN_10505 & _GEN_9838 ? io_writedata : CacheMem_2_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1885 = _GEN_10505 & _GEN_9842 ? io_writedata : CacheMem_2_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1886 = _GEN_10505 & _GEN_9846 ? io_writedata : CacheMem_2_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1887 = _GEN_10505 & _GEN_9850 ? io_writedata : CacheMem_2_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1888 = _GEN_10505 & _GEN_9854 ? io_writedata : CacheMem_2_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1889 = _GEN_10505 & _GEN_9858 ? io_writedata : CacheMem_2_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1890 = _GEN_10505 & _GEN_9862 ? io_writedata : CacheMem_2_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1891 = _GEN_10537 & _GEN_9866 ? io_writedata : CacheMem_2_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1892 = _GEN_10537 & _GEN_9838 ? io_writedata : CacheMem_2_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1893 = _GEN_10537 & _GEN_9842 ? io_writedata : CacheMem_2_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1894 = _GEN_10537 & _GEN_9846 ? io_writedata : CacheMem_2_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1895 = _GEN_10537 & _GEN_9850 ? io_writedata : CacheMem_2_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1896 = _GEN_10537 & _GEN_9854 ? io_writedata : CacheMem_2_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1897 = _GEN_10537 & _GEN_9858 ? io_writedata : CacheMem_2_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1898 = _GEN_10537 & _GEN_9862 ? io_writedata : CacheMem_2_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1899 = _GEN_10569 & _GEN_9866 ? io_writedata : CacheMem_2_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1900 = _GEN_10569 & _GEN_9838 ? io_writedata : CacheMem_2_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1901 = _GEN_10569 & _GEN_9842 ? io_writedata : CacheMem_2_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1902 = _GEN_10569 & _GEN_9846 ? io_writedata : CacheMem_2_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1903 = _GEN_10569 & _GEN_9850 ? io_writedata : CacheMem_2_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1904 = _GEN_10569 & _GEN_9854 ? io_writedata : CacheMem_2_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1905 = _GEN_10569 & _GEN_9858 ? io_writedata : CacheMem_2_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1906 = _GEN_10569 & _GEN_9862 ? io_writedata : CacheMem_2_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1907 = _GEN_10601 & _GEN_9866 ? io_writedata : CacheMem_3_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1908 = _GEN_10601 & _GEN_9838 ? io_writedata : CacheMem_3_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1909 = _GEN_10601 & _GEN_9842 ? io_writedata : CacheMem_3_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1910 = _GEN_10601 & _GEN_9846 ? io_writedata : CacheMem_3_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1911 = _GEN_10601 & _GEN_9850 ? io_writedata : CacheMem_3_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1912 = _GEN_10601 & _GEN_9854 ? io_writedata : CacheMem_3_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1913 = _GEN_10601 & _GEN_9858 ? io_writedata : CacheMem_3_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1914 = _GEN_10601 & _GEN_9862 ? io_writedata : CacheMem_3_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1915 = _GEN_10633 & _GEN_9866 ? io_writedata : CacheMem_3_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1916 = _GEN_10633 & _GEN_9838 ? io_writedata : CacheMem_3_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1917 = _GEN_10633 & _GEN_9842 ? io_writedata : CacheMem_3_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1918 = _GEN_10633 & _GEN_9846 ? io_writedata : CacheMem_3_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1919 = _GEN_10633 & _GEN_9850 ? io_writedata : CacheMem_3_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1920 = _GEN_10633 & _GEN_9854 ? io_writedata : CacheMem_3_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1921 = _GEN_10633 & _GEN_9858 ? io_writedata : CacheMem_3_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1922 = _GEN_10633 & _GEN_9862 ? io_writedata : CacheMem_3_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1923 = _GEN_10665 & _GEN_9866 ? io_writedata : CacheMem_3_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1924 = _GEN_10665 & _GEN_9838 ? io_writedata : CacheMem_3_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1925 = _GEN_10665 & _GEN_9842 ? io_writedata : CacheMem_3_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1926 = _GEN_10665 & _GEN_9846 ? io_writedata : CacheMem_3_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1927 = _GEN_10665 & _GEN_9850 ? io_writedata : CacheMem_3_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1928 = _GEN_10665 & _GEN_9854 ? io_writedata : CacheMem_3_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1929 = _GEN_10665 & _GEN_9858 ? io_writedata : CacheMem_3_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1930 = _GEN_10665 & _GEN_9862 ? io_writedata : CacheMem_3_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1931 = _GEN_10697 & _GEN_9866 ? io_writedata : CacheMem_3_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1932 = _GEN_10697 & _GEN_9838 ? io_writedata : CacheMem_3_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1933 = _GEN_10697 & _GEN_9842 ? io_writedata : CacheMem_3_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1934 = _GEN_10697 & _GEN_9846 ? io_writedata : CacheMem_3_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1935 = _GEN_10697 & _GEN_9850 ? io_writedata : CacheMem_3_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1936 = _GEN_10697 & _GEN_9854 ? io_writedata : CacheMem_3_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1937 = _GEN_10697 & _GEN_9858 ? io_writedata : CacheMem_3_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1938 = _GEN_10697 & _GEN_9862 ? io_writedata : CacheMem_3_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1939 = _GEN_10729 & _GEN_9866 ? io_writedata : CacheMem_3_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1940 = _GEN_10729 & _GEN_9838 ? io_writedata : CacheMem_3_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1941 = _GEN_10729 & _GEN_9842 ? io_writedata : CacheMem_3_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1942 = _GEN_10729 & _GEN_9846 ? io_writedata : CacheMem_3_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1943 = _GEN_10729 & _GEN_9850 ? io_writedata : CacheMem_3_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1944 = _GEN_10729 & _GEN_9854 ? io_writedata : CacheMem_3_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1945 = _GEN_10729 & _GEN_9858 ? io_writedata : CacheMem_3_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1946 = _GEN_10729 & _GEN_9862 ? io_writedata : CacheMem_3_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1947 = _GEN_10761 & _GEN_9866 ? io_writedata : CacheMem_3_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1948 = _GEN_10761 & _GEN_9838 ? io_writedata : CacheMem_3_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1949 = _GEN_10761 & _GEN_9842 ? io_writedata : CacheMem_3_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1950 = _GEN_10761 & _GEN_9846 ? io_writedata : CacheMem_3_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1951 = _GEN_10761 & _GEN_9850 ? io_writedata : CacheMem_3_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1952 = _GEN_10761 & _GEN_9854 ? io_writedata : CacheMem_3_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1953 = _GEN_10761 & _GEN_9858 ? io_writedata : CacheMem_3_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1954 = _GEN_10761 & _GEN_9862 ? io_writedata : CacheMem_3_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1955 = _GEN_10793 & _GEN_9866 ? io_writedata : CacheMem_3_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1956 = _GEN_10793 & _GEN_9838 ? io_writedata : CacheMem_3_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1957 = _GEN_10793 & _GEN_9842 ? io_writedata : CacheMem_3_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1958 = _GEN_10793 & _GEN_9846 ? io_writedata : CacheMem_3_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1959 = _GEN_10793 & _GEN_9850 ? io_writedata : CacheMem_3_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1960 = _GEN_10793 & _GEN_9854 ? io_writedata : CacheMem_3_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1961 = _GEN_10793 & _GEN_9858 ? io_writedata : CacheMem_3_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1962 = _GEN_10793 & _GEN_9862 ? io_writedata : CacheMem_3_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1963 = _GEN_10825 & _GEN_9866 ? io_writedata : CacheMem_3_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1964 = _GEN_10825 & _GEN_9838 ? io_writedata : CacheMem_3_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1965 = _GEN_10825 & _GEN_9842 ? io_writedata : CacheMem_3_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1966 = _GEN_10825 & _GEN_9846 ? io_writedata : CacheMem_3_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1967 = _GEN_10825 & _GEN_9850 ? io_writedata : CacheMem_3_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1968 = _GEN_10825 & _GEN_9854 ? io_writedata : CacheMem_3_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1969 = _GEN_10825 & _GEN_9858 ? io_writedata : CacheMem_3_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1970 = _GEN_10825 & _GEN_9862 ? io_writedata : CacheMem_3_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1971 = _GEN_10857 & _GEN_9866 ? io_writedata : CacheMem_4_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1972 = _GEN_10857 & _GEN_9838 ? io_writedata : CacheMem_4_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1973 = _GEN_10857 & _GEN_9842 ? io_writedata : CacheMem_4_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1974 = _GEN_10857 & _GEN_9846 ? io_writedata : CacheMem_4_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1975 = _GEN_10857 & _GEN_9850 ? io_writedata : CacheMem_4_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1976 = _GEN_10857 & _GEN_9854 ? io_writedata : CacheMem_4_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1977 = _GEN_10857 & _GEN_9858 ? io_writedata : CacheMem_4_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1978 = _GEN_10857 & _GEN_9862 ? io_writedata : CacheMem_4_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1979 = _GEN_10889 & _GEN_9866 ? io_writedata : CacheMem_4_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1980 = _GEN_10889 & _GEN_9838 ? io_writedata : CacheMem_4_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1981 = _GEN_10889 & _GEN_9842 ? io_writedata : CacheMem_4_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1982 = _GEN_10889 & _GEN_9846 ? io_writedata : CacheMem_4_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1983 = _GEN_10889 & _GEN_9850 ? io_writedata : CacheMem_4_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1984 = _GEN_10889 & _GEN_9854 ? io_writedata : CacheMem_4_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1985 = _GEN_10889 & _GEN_9858 ? io_writedata : CacheMem_4_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1986 = _GEN_10889 & _GEN_9862 ? io_writedata : CacheMem_4_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1987 = _GEN_10921 & _GEN_9866 ? io_writedata : CacheMem_4_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1988 = _GEN_10921 & _GEN_9838 ? io_writedata : CacheMem_4_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1989 = _GEN_10921 & _GEN_9842 ? io_writedata : CacheMem_4_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1990 = _GEN_10921 & _GEN_9846 ? io_writedata : CacheMem_4_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1991 = _GEN_10921 & _GEN_9850 ? io_writedata : CacheMem_4_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1992 = _GEN_10921 & _GEN_9854 ? io_writedata : CacheMem_4_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1993 = _GEN_10921 & _GEN_9858 ? io_writedata : CacheMem_4_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1994 = _GEN_10921 & _GEN_9862 ? io_writedata : CacheMem_4_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1995 = _GEN_10953 & _GEN_9866 ? io_writedata : CacheMem_4_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1996 = _GEN_10953 & _GEN_9838 ? io_writedata : CacheMem_4_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1997 = _GEN_10953 & _GEN_9842 ? io_writedata : CacheMem_4_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1998 = _GEN_10953 & _GEN_9846 ? io_writedata : CacheMem_4_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_1999 = _GEN_10953 & _GEN_9850 ? io_writedata : CacheMem_4_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2000 = _GEN_10953 & _GEN_9854 ? io_writedata : CacheMem_4_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2001 = _GEN_10953 & _GEN_9858 ? io_writedata : CacheMem_4_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2002 = _GEN_10953 & _GEN_9862 ? io_writedata : CacheMem_4_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2003 = _GEN_10985 & _GEN_9866 ? io_writedata : CacheMem_4_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2004 = _GEN_10985 & _GEN_9838 ? io_writedata : CacheMem_4_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2005 = _GEN_10985 & _GEN_9842 ? io_writedata : CacheMem_4_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2006 = _GEN_10985 & _GEN_9846 ? io_writedata : CacheMem_4_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2007 = _GEN_10985 & _GEN_9850 ? io_writedata : CacheMem_4_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2008 = _GEN_10985 & _GEN_9854 ? io_writedata : CacheMem_4_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2009 = _GEN_10985 & _GEN_9858 ? io_writedata : CacheMem_4_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2010 = _GEN_10985 & _GEN_9862 ? io_writedata : CacheMem_4_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2011 = _GEN_11017 & _GEN_9866 ? io_writedata : CacheMem_4_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2012 = _GEN_11017 & _GEN_9838 ? io_writedata : CacheMem_4_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2013 = _GEN_11017 & _GEN_9842 ? io_writedata : CacheMem_4_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2014 = _GEN_11017 & _GEN_9846 ? io_writedata : CacheMem_4_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2015 = _GEN_11017 & _GEN_9850 ? io_writedata : CacheMem_4_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2016 = _GEN_11017 & _GEN_9854 ? io_writedata : CacheMem_4_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2017 = _GEN_11017 & _GEN_9858 ? io_writedata : CacheMem_4_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2018 = _GEN_11017 & _GEN_9862 ? io_writedata : CacheMem_4_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2019 = _GEN_11049 & _GEN_9866 ? io_writedata : CacheMem_4_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2020 = _GEN_11049 & _GEN_9838 ? io_writedata : CacheMem_4_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2021 = _GEN_11049 & _GEN_9842 ? io_writedata : CacheMem_4_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2022 = _GEN_11049 & _GEN_9846 ? io_writedata : CacheMem_4_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2023 = _GEN_11049 & _GEN_9850 ? io_writedata : CacheMem_4_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2024 = _GEN_11049 & _GEN_9854 ? io_writedata : CacheMem_4_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2025 = _GEN_11049 & _GEN_9858 ? io_writedata : CacheMem_4_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2026 = _GEN_11049 & _GEN_9862 ? io_writedata : CacheMem_4_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2027 = _GEN_11081 & _GEN_9866 ? io_writedata : CacheMem_4_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2028 = _GEN_11081 & _GEN_9838 ? io_writedata : CacheMem_4_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2029 = _GEN_11081 & _GEN_9842 ? io_writedata : CacheMem_4_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2030 = _GEN_11081 & _GEN_9846 ? io_writedata : CacheMem_4_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2031 = _GEN_11081 & _GEN_9850 ? io_writedata : CacheMem_4_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2032 = _GEN_11081 & _GEN_9854 ? io_writedata : CacheMem_4_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2033 = _GEN_11081 & _GEN_9858 ? io_writedata : CacheMem_4_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2034 = _GEN_11081 & _GEN_9862 ? io_writedata : CacheMem_4_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2035 = _GEN_11113 & _GEN_9866 ? io_writedata : CacheMem_5_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2036 = _GEN_11113 & _GEN_9838 ? io_writedata : CacheMem_5_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2037 = _GEN_11113 & _GEN_9842 ? io_writedata : CacheMem_5_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2038 = _GEN_11113 & _GEN_9846 ? io_writedata : CacheMem_5_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2039 = _GEN_11113 & _GEN_9850 ? io_writedata : CacheMem_5_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2040 = _GEN_11113 & _GEN_9854 ? io_writedata : CacheMem_5_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2041 = _GEN_11113 & _GEN_9858 ? io_writedata : CacheMem_5_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2042 = _GEN_11113 & _GEN_9862 ? io_writedata : CacheMem_5_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2043 = _GEN_11145 & _GEN_9866 ? io_writedata : CacheMem_5_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2044 = _GEN_11145 & _GEN_9838 ? io_writedata : CacheMem_5_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2045 = _GEN_11145 & _GEN_9842 ? io_writedata : CacheMem_5_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2046 = _GEN_11145 & _GEN_9846 ? io_writedata : CacheMem_5_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2047 = _GEN_11145 & _GEN_9850 ? io_writedata : CacheMem_5_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2048 = _GEN_11145 & _GEN_9854 ? io_writedata : CacheMem_5_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2049 = _GEN_11145 & _GEN_9858 ? io_writedata : CacheMem_5_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2050 = _GEN_11145 & _GEN_9862 ? io_writedata : CacheMem_5_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2051 = _GEN_11177 & _GEN_9866 ? io_writedata : CacheMem_5_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2052 = _GEN_11177 & _GEN_9838 ? io_writedata : CacheMem_5_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2053 = _GEN_11177 & _GEN_9842 ? io_writedata : CacheMem_5_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2054 = _GEN_11177 & _GEN_9846 ? io_writedata : CacheMem_5_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2055 = _GEN_11177 & _GEN_9850 ? io_writedata : CacheMem_5_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2056 = _GEN_11177 & _GEN_9854 ? io_writedata : CacheMem_5_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2057 = _GEN_11177 & _GEN_9858 ? io_writedata : CacheMem_5_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2058 = _GEN_11177 & _GEN_9862 ? io_writedata : CacheMem_5_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2059 = _GEN_11209 & _GEN_9866 ? io_writedata : CacheMem_5_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2060 = _GEN_11209 & _GEN_9838 ? io_writedata : CacheMem_5_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2061 = _GEN_11209 & _GEN_9842 ? io_writedata : CacheMem_5_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2062 = _GEN_11209 & _GEN_9846 ? io_writedata : CacheMem_5_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2063 = _GEN_11209 & _GEN_9850 ? io_writedata : CacheMem_5_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2064 = _GEN_11209 & _GEN_9854 ? io_writedata : CacheMem_5_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2065 = _GEN_11209 & _GEN_9858 ? io_writedata : CacheMem_5_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2066 = _GEN_11209 & _GEN_9862 ? io_writedata : CacheMem_5_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2067 = _GEN_11241 & _GEN_9866 ? io_writedata : CacheMem_5_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2068 = _GEN_11241 & _GEN_9838 ? io_writedata : CacheMem_5_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2069 = _GEN_11241 & _GEN_9842 ? io_writedata : CacheMem_5_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2070 = _GEN_11241 & _GEN_9846 ? io_writedata : CacheMem_5_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2071 = _GEN_11241 & _GEN_9850 ? io_writedata : CacheMem_5_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2072 = _GEN_11241 & _GEN_9854 ? io_writedata : CacheMem_5_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2073 = _GEN_11241 & _GEN_9858 ? io_writedata : CacheMem_5_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2074 = _GEN_11241 & _GEN_9862 ? io_writedata : CacheMem_5_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2075 = _GEN_11273 & _GEN_9866 ? io_writedata : CacheMem_5_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2076 = _GEN_11273 & _GEN_9838 ? io_writedata : CacheMem_5_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2077 = _GEN_11273 & _GEN_9842 ? io_writedata : CacheMem_5_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2078 = _GEN_11273 & _GEN_9846 ? io_writedata : CacheMem_5_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2079 = _GEN_11273 & _GEN_9850 ? io_writedata : CacheMem_5_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2080 = _GEN_11273 & _GEN_9854 ? io_writedata : CacheMem_5_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2081 = _GEN_11273 & _GEN_9858 ? io_writedata : CacheMem_5_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2082 = _GEN_11273 & _GEN_9862 ? io_writedata : CacheMem_5_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2083 = _GEN_11305 & _GEN_9866 ? io_writedata : CacheMem_5_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2084 = _GEN_11305 & _GEN_9838 ? io_writedata : CacheMem_5_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2085 = _GEN_11305 & _GEN_9842 ? io_writedata : CacheMem_5_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2086 = _GEN_11305 & _GEN_9846 ? io_writedata : CacheMem_5_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2087 = _GEN_11305 & _GEN_9850 ? io_writedata : CacheMem_5_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2088 = _GEN_11305 & _GEN_9854 ? io_writedata : CacheMem_5_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2089 = _GEN_11305 & _GEN_9858 ? io_writedata : CacheMem_5_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2090 = _GEN_11305 & _GEN_9862 ? io_writedata : CacheMem_5_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2091 = _GEN_11337 & _GEN_9866 ? io_writedata : CacheMem_5_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2092 = _GEN_11337 & _GEN_9838 ? io_writedata : CacheMem_5_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2093 = _GEN_11337 & _GEN_9842 ? io_writedata : CacheMem_5_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2094 = _GEN_11337 & _GEN_9846 ? io_writedata : CacheMem_5_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2095 = _GEN_11337 & _GEN_9850 ? io_writedata : CacheMem_5_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2096 = _GEN_11337 & _GEN_9854 ? io_writedata : CacheMem_5_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2097 = _GEN_11337 & _GEN_9858 ? io_writedata : CacheMem_5_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2098 = _GEN_11337 & _GEN_9862 ? io_writedata : CacheMem_5_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2099 = _GEN_11369 & _GEN_9866 ? io_writedata : CacheMem_6_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2100 = _GEN_11369 & _GEN_9838 ? io_writedata : CacheMem_6_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2101 = _GEN_11369 & _GEN_9842 ? io_writedata : CacheMem_6_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2102 = _GEN_11369 & _GEN_9846 ? io_writedata : CacheMem_6_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2103 = _GEN_11369 & _GEN_9850 ? io_writedata : CacheMem_6_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2104 = _GEN_11369 & _GEN_9854 ? io_writedata : CacheMem_6_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2105 = _GEN_11369 & _GEN_9858 ? io_writedata : CacheMem_6_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2106 = _GEN_11369 & _GEN_9862 ? io_writedata : CacheMem_6_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2107 = _GEN_11401 & _GEN_9866 ? io_writedata : CacheMem_6_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2108 = _GEN_11401 & _GEN_9838 ? io_writedata : CacheMem_6_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2109 = _GEN_11401 & _GEN_9842 ? io_writedata : CacheMem_6_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2110 = _GEN_11401 & _GEN_9846 ? io_writedata : CacheMem_6_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2111 = _GEN_11401 & _GEN_9850 ? io_writedata : CacheMem_6_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2112 = _GEN_11401 & _GEN_9854 ? io_writedata : CacheMem_6_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2113 = _GEN_11401 & _GEN_9858 ? io_writedata : CacheMem_6_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2114 = _GEN_11401 & _GEN_9862 ? io_writedata : CacheMem_6_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2115 = _GEN_11433 & _GEN_9866 ? io_writedata : CacheMem_6_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2116 = _GEN_11433 & _GEN_9838 ? io_writedata : CacheMem_6_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2117 = _GEN_11433 & _GEN_9842 ? io_writedata : CacheMem_6_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2118 = _GEN_11433 & _GEN_9846 ? io_writedata : CacheMem_6_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2119 = _GEN_11433 & _GEN_9850 ? io_writedata : CacheMem_6_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2120 = _GEN_11433 & _GEN_9854 ? io_writedata : CacheMem_6_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2121 = _GEN_11433 & _GEN_9858 ? io_writedata : CacheMem_6_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2122 = _GEN_11433 & _GEN_9862 ? io_writedata : CacheMem_6_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2123 = _GEN_11465 & _GEN_9866 ? io_writedata : CacheMem_6_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2124 = _GEN_11465 & _GEN_9838 ? io_writedata : CacheMem_6_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2125 = _GEN_11465 & _GEN_9842 ? io_writedata : CacheMem_6_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2126 = _GEN_11465 & _GEN_9846 ? io_writedata : CacheMem_6_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2127 = _GEN_11465 & _GEN_9850 ? io_writedata : CacheMem_6_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2128 = _GEN_11465 & _GEN_9854 ? io_writedata : CacheMem_6_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2129 = _GEN_11465 & _GEN_9858 ? io_writedata : CacheMem_6_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2130 = _GEN_11465 & _GEN_9862 ? io_writedata : CacheMem_6_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2131 = _GEN_11497 & _GEN_9866 ? io_writedata : CacheMem_6_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2132 = _GEN_11497 & _GEN_9838 ? io_writedata : CacheMem_6_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2133 = _GEN_11497 & _GEN_9842 ? io_writedata : CacheMem_6_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2134 = _GEN_11497 & _GEN_9846 ? io_writedata : CacheMem_6_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2135 = _GEN_11497 & _GEN_9850 ? io_writedata : CacheMem_6_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2136 = _GEN_11497 & _GEN_9854 ? io_writedata : CacheMem_6_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2137 = _GEN_11497 & _GEN_9858 ? io_writedata : CacheMem_6_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2138 = _GEN_11497 & _GEN_9862 ? io_writedata : CacheMem_6_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2139 = _GEN_11529 & _GEN_9866 ? io_writedata : CacheMem_6_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2140 = _GEN_11529 & _GEN_9838 ? io_writedata : CacheMem_6_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2141 = _GEN_11529 & _GEN_9842 ? io_writedata : CacheMem_6_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2142 = _GEN_11529 & _GEN_9846 ? io_writedata : CacheMem_6_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2143 = _GEN_11529 & _GEN_9850 ? io_writedata : CacheMem_6_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2144 = _GEN_11529 & _GEN_9854 ? io_writedata : CacheMem_6_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2145 = _GEN_11529 & _GEN_9858 ? io_writedata : CacheMem_6_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2146 = _GEN_11529 & _GEN_9862 ? io_writedata : CacheMem_6_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2147 = _GEN_11561 & _GEN_9866 ? io_writedata : CacheMem_6_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2148 = _GEN_11561 & _GEN_9838 ? io_writedata : CacheMem_6_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2149 = _GEN_11561 & _GEN_9842 ? io_writedata : CacheMem_6_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2150 = _GEN_11561 & _GEN_9846 ? io_writedata : CacheMem_6_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2151 = _GEN_11561 & _GEN_9850 ? io_writedata : CacheMem_6_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2152 = _GEN_11561 & _GEN_9854 ? io_writedata : CacheMem_6_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2153 = _GEN_11561 & _GEN_9858 ? io_writedata : CacheMem_6_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2154 = _GEN_11561 & _GEN_9862 ? io_writedata : CacheMem_6_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2155 = _GEN_11593 & _GEN_9866 ? io_writedata : CacheMem_6_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2156 = _GEN_11593 & _GEN_9838 ? io_writedata : CacheMem_6_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2157 = _GEN_11593 & _GEN_9842 ? io_writedata : CacheMem_6_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2158 = _GEN_11593 & _GEN_9846 ? io_writedata : CacheMem_6_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2159 = _GEN_11593 & _GEN_9850 ? io_writedata : CacheMem_6_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2160 = _GEN_11593 & _GEN_9854 ? io_writedata : CacheMem_6_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2161 = _GEN_11593 & _GEN_9858 ? io_writedata : CacheMem_6_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2162 = _GEN_11593 & _GEN_9862 ? io_writedata : CacheMem_6_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2163 = _GEN_11625 & _GEN_9866 ? io_writedata : CacheMem_7_0_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2164 = _GEN_11625 & _GEN_9838 ? io_writedata : CacheMem_7_0_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2165 = _GEN_11625 & _GEN_9842 ? io_writedata : CacheMem_7_0_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2166 = _GEN_11625 & _GEN_9846 ? io_writedata : CacheMem_7_0_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2167 = _GEN_11625 & _GEN_9850 ? io_writedata : CacheMem_7_0_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2168 = _GEN_11625 & _GEN_9854 ? io_writedata : CacheMem_7_0_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2169 = _GEN_11625 & _GEN_9858 ? io_writedata : CacheMem_7_0_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2170 = _GEN_11625 & _GEN_9862 ? io_writedata : CacheMem_7_0_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2171 = _GEN_11657 & _GEN_9866 ? io_writedata : CacheMem_7_1_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2172 = _GEN_11657 & _GEN_9838 ? io_writedata : CacheMem_7_1_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2173 = _GEN_11657 & _GEN_9842 ? io_writedata : CacheMem_7_1_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2174 = _GEN_11657 & _GEN_9846 ? io_writedata : CacheMem_7_1_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2175 = _GEN_11657 & _GEN_9850 ? io_writedata : CacheMem_7_1_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2176 = _GEN_11657 & _GEN_9854 ? io_writedata : CacheMem_7_1_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2177 = _GEN_11657 & _GEN_9858 ? io_writedata : CacheMem_7_1_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2178 = _GEN_11657 & _GEN_9862 ? io_writedata : CacheMem_7_1_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2179 = _GEN_11689 & _GEN_9866 ? io_writedata : CacheMem_7_2_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2180 = _GEN_11689 & _GEN_9838 ? io_writedata : CacheMem_7_2_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2181 = _GEN_11689 & _GEN_9842 ? io_writedata : CacheMem_7_2_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2182 = _GEN_11689 & _GEN_9846 ? io_writedata : CacheMem_7_2_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2183 = _GEN_11689 & _GEN_9850 ? io_writedata : CacheMem_7_2_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2184 = _GEN_11689 & _GEN_9854 ? io_writedata : CacheMem_7_2_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2185 = _GEN_11689 & _GEN_9858 ? io_writedata : CacheMem_7_2_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2186 = _GEN_11689 & _GEN_9862 ? io_writedata : CacheMem_7_2_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2187 = _GEN_11721 & _GEN_9866 ? io_writedata : CacheMem_7_3_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2188 = _GEN_11721 & _GEN_9838 ? io_writedata : CacheMem_7_3_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2189 = _GEN_11721 & _GEN_9842 ? io_writedata : CacheMem_7_3_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2190 = _GEN_11721 & _GEN_9846 ? io_writedata : CacheMem_7_3_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2191 = _GEN_11721 & _GEN_9850 ? io_writedata : CacheMem_7_3_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2192 = _GEN_11721 & _GEN_9854 ? io_writedata : CacheMem_7_3_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2193 = _GEN_11721 & _GEN_9858 ? io_writedata : CacheMem_7_3_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2194 = _GEN_11721 & _GEN_9862 ? io_writedata : CacheMem_7_3_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2195 = _GEN_11753 & _GEN_9866 ? io_writedata : CacheMem_7_4_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2196 = _GEN_11753 & _GEN_9838 ? io_writedata : CacheMem_7_4_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2197 = _GEN_11753 & _GEN_9842 ? io_writedata : CacheMem_7_4_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2198 = _GEN_11753 & _GEN_9846 ? io_writedata : CacheMem_7_4_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2199 = _GEN_11753 & _GEN_9850 ? io_writedata : CacheMem_7_4_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2200 = _GEN_11753 & _GEN_9854 ? io_writedata : CacheMem_7_4_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2201 = _GEN_11753 & _GEN_9858 ? io_writedata : CacheMem_7_4_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2202 = _GEN_11753 & _GEN_9862 ? io_writedata : CacheMem_7_4_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2203 = _GEN_11785 & _GEN_9866 ? io_writedata : CacheMem_7_5_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2204 = _GEN_11785 & _GEN_9838 ? io_writedata : CacheMem_7_5_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2205 = _GEN_11785 & _GEN_9842 ? io_writedata : CacheMem_7_5_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2206 = _GEN_11785 & _GEN_9846 ? io_writedata : CacheMem_7_5_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2207 = _GEN_11785 & _GEN_9850 ? io_writedata : CacheMem_7_5_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2208 = _GEN_11785 & _GEN_9854 ? io_writedata : CacheMem_7_5_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2209 = _GEN_11785 & _GEN_9858 ? io_writedata : CacheMem_7_5_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2210 = _GEN_11785 & _GEN_9862 ? io_writedata : CacheMem_7_5_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2211 = _GEN_11817 & _GEN_9866 ? io_writedata : CacheMem_7_6_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2212 = _GEN_11817 & _GEN_9838 ? io_writedata : CacheMem_7_6_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2213 = _GEN_11817 & _GEN_9842 ? io_writedata : CacheMem_7_6_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2214 = _GEN_11817 & _GEN_9846 ? io_writedata : CacheMem_7_6_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2215 = _GEN_11817 & _GEN_9850 ? io_writedata : CacheMem_7_6_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2216 = _GEN_11817 & _GEN_9854 ? io_writedata : CacheMem_7_6_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2217 = _GEN_11817 & _GEN_9858 ? io_writedata : CacheMem_7_6_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2218 = _GEN_11817 & _GEN_9862 ? io_writedata : CacheMem_7_6_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2219 = _GEN_11849 & _GEN_9866 ? io_writedata : CacheMem_7_7_0; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2220 = _GEN_11849 & _GEN_9838 ? io_writedata : CacheMem_7_7_1; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2221 = _GEN_11849 & _GEN_9842 ? io_writedata : CacheMem_7_7_2; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2222 = _GEN_11849 & _GEN_9846 ? io_writedata : CacheMem_7_7_3; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2223 = _GEN_11849 & _GEN_9850 ? io_writedata : CacheMem_7_7_4; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2224 = _GEN_11849 & _GEN_9854 ? io_writedata : CacheMem_7_7_5; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2225 = _GEN_11849 & _GEN_9858 ? io_writedata : CacheMem_7_7_6; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2226 = _GEN_11849 & _GEN_9862 ? io_writedata : CacheMem_7_7_7; // @[Cache.scala 141:{54,54} 53:25]
  wire [31:0] _GEN_2227 = 4'hf == io_writeMask ? _GEN_1715 : CacheMem_0_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2228 = 4'hf == io_writeMask ? _GEN_1716 : CacheMem_0_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2229 = 4'hf == io_writeMask ? _GEN_1717 : CacheMem_0_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2230 = 4'hf == io_writeMask ? _GEN_1718 : CacheMem_0_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2231 = 4'hf == io_writeMask ? _GEN_1719 : CacheMem_0_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2232 = 4'hf == io_writeMask ? _GEN_1720 : CacheMem_0_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2233 = 4'hf == io_writeMask ? _GEN_1721 : CacheMem_0_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2234 = 4'hf == io_writeMask ? _GEN_1722 : CacheMem_0_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2235 = 4'hf == io_writeMask ? _GEN_1723 : CacheMem_0_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2236 = 4'hf == io_writeMask ? _GEN_1724 : CacheMem_0_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2237 = 4'hf == io_writeMask ? _GEN_1725 : CacheMem_0_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2238 = 4'hf == io_writeMask ? _GEN_1726 : CacheMem_0_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2239 = 4'hf == io_writeMask ? _GEN_1727 : CacheMem_0_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2240 = 4'hf == io_writeMask ? _GEN_1728 : CacheMem_0_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2241 = 4'hf == io_writeMask ? _GEN_1729 : CacheMem_0_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2242 = 4'hf == io_writeMask ? _GEN_1730 : CacheMem_0_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2243 = 4'hf == io_writeMask ? _GEN_1731 : CacheMem_0_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2244 = 4'hf == io_writeMask ? _GEN_1732 : CacheMem_0_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2245 = 4'hf == io_writeMask ? _GEN_1733 : CacheMem_0_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2246 = 4'hf == io_writeMask ? _GEN_1734 : CacheMem_0_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2247 = 4'hf == io_writeMask ? _GEN_1735 : CacheMem_0_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2248 = 4'hf == io_writeMask ? _GEN_1736 : CacheMem_0_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2249 = 4'hf == io_writeMask ? _GEN_1737 : CacheMem_0_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2250 = 4'hf == io_writeMask ? _GEN_1738 : CacheMem_0_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2251 = 4'hf == io_writeMask ? _GEN_1739 : CacheMem_0_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2252 = 4'hf == io_writeMask ? _GEN_1740 : CacheMem_0_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2253 = 4'hf == io_writeMask ? _GEN_1741 : CacheMem_0_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2254 = 4'hf == io_writeMask ? _GEN_1742 : CacheMem_0_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2255 = 4'hf == io_writeMask ? _GEN_1743 : CacheMem_0_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2256 = 4'hf == io_writeMask ? _GEN_1744 : CacheMem_0_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2257 = 4'hf == io_writeMask ? _GEN_1745 : CacheMem_0_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2258 = 4'hf == io_writeMask ? _GEN_1746 : CacheMem_0_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2259 = 4'hf == io_writeMask ? _GEN_1747 : CacheMem_0_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2260 = 4'hf == io_writeMask ? _GEN_1748 : CacheMem_0_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2261 = 4'hf == io_writeMask ? _GEN_1749 : CacheMem_0_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2262 = 4'hf == io_writeMask ? _GEN_1750 : CacheMem_0_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2263 = 4'hf == io_writeMask ? _GEN_1751 : CacheMem_0_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2264 = 4'hf == io_writeMask ? _GEN_1752 : CacheMem_0_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2265 = 4'hf == io_writeMask ? _GEN_1753 : CacheMem_0_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2266 = 4'hf == io_writeMask ? _GEN_1754 : CacheMem_0_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2267 = 4'hf == io_writeMask ? _GEN_1755 : CacheMem_0_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2268 = 4'hf == io_writeMask ? _GEN_1756 : CacheMem_0_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2269 = 4'hf == io_writeMask ? _GEN_1757 : CacheMem_0_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2270 = 4'hf == io_writeMask ? _GEN_1758 : CacheMem_0_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2271 = 4'hf == io_writeMask ? _GEN_1759 : CacheMem_0_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2272 = 4'hf == io_writeMask ? _GEN_1760 : CacheMem_0_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2273 = 4'hf == io_writeMask ? _GEN_1761 : CacheMem_0_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2274 = 4'hf == io_writeMask ? _GEN_1762 : CacheMem_0_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2275 = 4'hf == io_writeMask ? _GEN_1763 : CacheMem_0_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2276 = 4'hf == io_writeMask ? _GEN_1764 : CacheMem_0_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2277 = 4'hf == io_writeMask ? _GEN_1765 : CacheMem_0_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2278 = 4'hf == io_writeMask ? _GEN_1766 : CacheMem_0_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2279 = 4'hf == io_writeMask ? _GEN_1767 : CacheMem_0_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2280 = 4'hf == io_writeMask ? _GEN_1768 : CacheMem_0_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2281 = 4'hf == io_writeMask ? _GEN_1769 : CacheMem_0_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2282 = 4'hf == io_writeMask ? _GEN_1770 : CacheMem_0_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2283 = 4'hf == io_writeMask ? _GEN_1771 : CacheMem_0_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2284 = 4'hf == io_writeMask ? _GEN_1772 : CacheMem_0_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2285 = 4'hf == io_writeMask ? _GEN_1773 : CacheMem_0_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2286 = 4'hf == io_writeMask ? _GEN_1774 : CacheMem_0_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2287 = 4'hf == io_writeMask ? _GEN_1775 : CacheMem_0_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2288 = 4'hf == io_writeMask ? _GEN_1776 : CacheMem_0_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2289 = 4'hf == io_writeMask ? _GEN_1777 : CacheMem_0_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2290 = 4'hf == io_writeMask ? _GEN_1778 : CacheMem_0_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2291 = 4'hf == io_writeMask ? _GEN_1779 : CacheMem_1_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2292 = 4'hf == io_writeMask ? _GEN_1780 : CacheMem_1_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2293 = 4'hf == io_writeMask ? _GEN_1781 : CacheMem_1_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2294 = 4'hf == io_writeMask ? _GEN_1782 : CacheMem_1_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2295 = 4'hf == io_writeMask ? _GEN_1783 : CacheMem_1_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2296 = 4'hf == io_writeMask ? _GEN_1784 : CacheMem_1_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2297 = 4'hf == io_writeMask ? _GEN_1785 : CacheMem_1_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2298 = 4'hf == io_writeMask ? _GEN_1786 : CacheMem_1_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2299 = 4'hf == io_writeMask ? _GEN_1787 : CacheMem_1_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2300 = 4'hf == io_writeMask ? _GEN_1788 : CacheMem_1_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2301 = 4'hf == io_writeMask ? _GEN_1789 : CacheMem_1_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2302 = 4'hf == io_writeMask ? _GEN_1790 : CacheMem_1_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2303 = 4'hf == io_writeMask ? _GEN_1791 : CacheMem_1_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2304 = 4'hf == io_writeMask ? _GEN_1792 : CacheMem_1_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2305 = 4'hf == io_writeMask ? _GEN_1793 : CacheMem_1_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2306 = 4'hf == io_writeMask ? _GEN_1794 : CacheMem_1_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2307 = 4'hf == io_writeMask ? _GEN_1795 : CacheMem_1_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2308 = 4'hf == io_writeMask ? _GEN_1796 : CacheMem_1_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2309 = 4'hf == io_writeMask ? _GEN_1797 : CacheMem_1_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2310 = 4'hf == io_writeMask ? _GEN_1798 : CacheMem_1_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2311 = 4'hf == io_writeMask ? _GEN_1799 : CacheMem_1_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2312 = 4'hf == io_writeMask ? _GEN_1800 : CacheMem_1_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2313 = 4'hf == io_writeMask ? _GEN_1801 : CacheMem_1_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2314 = 4'hf == io_writeMask ? _GEN_1802 : CacheMem_1_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2315 = 4'hf == io_writeMask ? _GEN_1803 : CacheMem_1_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2316 = 4'hf == io_writeMask ? _GEN_1804 : CacheMem_1_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2317 = 4'hf == io_writeMask ? _GEN_1805 : CacheMem_1_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2318 = 4'hf == io_writeMask ? _GEN_1806 : CacheMem_1_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2319 = 4'hf == io_writeMask ? _GEN_1807 : CacheMem_1_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2320 = 4'hf == io_writeMask ? _GEN_1808 : CacheMem_1_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2321 = 4'hf == io_writeMask ? _GEN_1809 : CacheMem_1_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2322 = 4'hf == io_writeMask ? _GEN_1810 : CacheMem_1_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2323 = 4'hf == io_writeMask ? _GEN_1811 : CacheMem_1_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2324 = 4'hf == io_writeMask ? _GEN_1812 : CacheMem_1_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2325 = 4'hf == io_writeMask ? _GEN_1813 : CacheMem_1_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2326 = 4'hf == io_writeMask ? _GEN_1814 : CacheMem_1_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2327 = 4'hf == io_writeMask ? _GEN_1815 : CacheMem_1_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2328 = 4'hf == io_writeMask ? _GEN_1816 : CacheMem_1_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2329 = 4'hf == io_writeMask ? _GEN_1817 : CacheMem_1_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2330 = 4'hf == io_writeMask ? _GEN_1818 : CacheMem_1_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2331 = 4'hf == io_writeMask ? _GEN_1819 : CacheMem_1_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2332 = 4'hf == io_writeMask ? _GEN_1820 : CacheMem_1_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2333 = 4'hf == io_writeMask ? _GEN_1821 : CacheMem_1_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2334 = 4'hf == io_writeMask ? _GEN_1822 : CacheMem_1_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2335 = 4'hf == io_writeMask ? _GEN_1823 : CacheMem_1_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2336 = 4'hf == io_writeMask ? _GEN_1824 : CacheMem_1_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2337 = 4'hf == io_writeMask ? _GEN_1825 : CacheMem_1_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2338 = 4'hf == io_writeMask ? _GEN_1826 : CacheMem_1_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2339 = 4'hf == io_writeMask ? _GEN_1827 : CacheMem_1_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2340 = 4'hf == io_writeMask ? _GEN_1828 : CacheMem_1_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2341 = 4'hf == io_writeMask ? _GEN_1829 : CacheMem_1_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2342 = 4'hf == io_writeMask ? _GEN_1830 : CacheMem_1_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2343 = 4'hf == io_writeMask ? _GEN_1831 : CacheMem_1_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2344 = 4'hf == io_writeMask ? _GEN_1832 : CacheMem_1_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2345 = 4'hf == io_writeMask ? _GEN_1833 : CacheMem_1_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2346 = 4'hf == io_writeMask ? _GEN_1834 : CacheMem_1_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2347 = 4'hf == io_writeMask ? _GEN_1835 : CacheMem_1_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2348 = 4'hf == io_writeMask ? _GEN_1836 : CacheMem_1_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2349 = 4'hf == io_writeMask ? _GEN_1837 : CacheMem_1_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2350 = 4'hf == io_writeMask ? _GEN_1838 : CacheMem_1_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2351 = 4'hf == io_writeMask ? _GEN_1839 : CacheMem_1_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2352 = 4'hf == io_writeMask ? _GEN_1840 : CacheMem_1_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2353 = 4'hf == io_writeMask ? _GEN_1841 : CacheMem_1_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2354 = 4'hf == io_writeMask ? _GEN_1842 : CacheMem_1_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2355 = 4'hf == io_writeMask ? _GEN_1843 : CacheMem_2_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2356 = 4'hf == io_writeMask ? _GEN_1844 : CacheMem_2_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2357 = 4'hf == io_writeMask ? _GEN_1845 : CacheMem_2_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2358 = 4'hf == io_writeMask ? _GEN_1846 : CacheMem_2_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2359 = 4'hf == io_writeMask ? _GEN_1847 : CacheMem_2_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2360 = 4'hf == io_writeMask ? _GEN_1848 : CacheMem_2_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2361 = 4'hf == io_writeMask ? _GEN_1849 : CacheMem_2_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2362 = 4'hf == io_writeMask ? _GEN_1850 : CacheMem_2_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2363 = 4'hf == io_writeMask ? _GEN_1851 : CacheMem_2_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2364 = 4'hf == io_writeMask ? _GEN_1852 : CacheMem_2_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2365 = 4'hf == io_writeMask ? _GEN_1853 : CacheMem_2_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2366 = 4'hf == io_writeMask ? _GEN_1854 : CacheMem_2_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2367 = 4'hf == io_writeMask ? _GEN_1855 : CacheMem_2_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2368 = 4'hf == io_writeMask ? _GEN_1856 : CacheMem_2_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2369 = 4'hf == io_writeMask ? _GEN_1857 : CacheMem_2_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2370 = 4'hf == io_writeMask ? _GEN_1858 : CacheMem_2_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2371 = 4'hf == io_writeMask ? _GEN_1859 : CacheMem_2_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2372 = 4'hf == io_writeMask ? _GEN_1860 : CacheMem_2_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2373 = 4'hf == io_writeMask ? _GEN_1861 : CacheMem_2_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2374 = 4'hf == io_writeMask ? _GEN_1862 : CacheMem_2_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2375 = 4'hf == io_writeMask ? _GEN_1863 : CacheMem_2_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2376 = 4'hf == io_writeMask ? _GEN_1864 : CacheMem_2_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2377 = 4'hf == io_writeMask ? _GEN_1865 : CacheMem_2_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2378 = 4'hf == io_writeMask ? _GEN_1866 : CacheMem_2_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2379 = 4'hf == io_writeMask ? _GEN_1867 : CacheMem_2_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2380 = 4'hf == io_writeMask ? _GEN_1868 : CacheMem_2_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2381 = 4'hf == io_writeMask ? _GEN_1869 : CacheMem_2_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2382 = 4'hf == io_writeMask ? _GEN_1870 : CacheMem_2_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2383 = 4'hf == io_writeMask ? _GEN_1871 : CacheMem_2_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2384 = 4'hf == io_writeMask ? _GEN_1872 : CacheMem_2_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2385 = 4'hf == io_writeMask ? _GEN_1873 : CacheMem_2_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2386 = 4'hf == io_writeMask ? _GEN_1874 : CacheMem_2_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2387 = 4'hf == io_writeMask ? _GEN_1875 : CacheMem_2_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2388 = 4'hf == io_writeMask ? _GEN_1876 : CacheMem_2_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2389 = 4'hf == io_writeMask ? _GEN_1877 : CacheMem_2_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2390 = 4'hf == io_writeMask ? _GEN_1878 : CacheMem_2_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2391 = 4'hf == io_writeMask ? _GEN_1879 : CacheMem_2_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2392 = 4'hf == io_writeMask ? _GEN_1880 : CacheMem_2_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2393 = 4'hf == io_writeMask ? _GEN_1881 : CacheMem_2_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2394 = 4'hf == io_writeMask ? _GEN_1882 : CacheMem_2_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2395 = 4'hf == io_writeMask ? _GEN_1883 : CacheMem_2_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2396 = 4'hf == io_writeMask ? _GEN_1884 : CacheMem_2_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2397 = 4'hf == io_writeMask ? _GEN_1885 : CacheMem_2_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2398 = 4'hf == io_writeMask ? _GEN_1886 : CacheMem_2_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2399 = 4'hf == io_writeMask ? _GEN_1887 : CacheMem_2_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2400 = 4'hf == io_writeMask ? _GEN_1888 : CacheMem_2_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2401 = 4'hf == io_writeMask ? _GEN_1889 : CacheMem_2_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2402 = 4'hf == io_writeMask ? _GEN_1890 : CacheMem_2_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2403 = 4'hf == io_writeMask ? _GEN_1891 : CacheMem_2_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2404 = 4'hf == io_writeMask ? _GEN_1892 : CacheMem_2_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2405 = 4'hf == io_writeMask ? _GEN_1893 : CacheMem_2_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2406 = 4'hf == io_writeMask ? _GEN_1894 : CacheMem_2_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2407 = 4'hf == io_writeMask ? _GEN_1895 : CacheMem_2_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2408 = 4'hf == io_writeMask ? _GEN_1896 : CacheMem_2_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2409 = 4'hf == io_writeMask ? _GEN_1897 : CacheMem_2_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2410 = 4'hf == io_writeMask ? _GEN_1898 : CacheMem_2_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2411 = 4'hf == io_writeMask ? _GEN_1899 : CacheMem_2_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2412 = 4'hf == io_writeMask ? _GEN_1900 : CacheMem_2_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2413 = 4'hf == io_writeMask ? _GEN_1901 : CacheMem_2_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2414 = 4'hf == io_writeMask ? _GEN_1902 : CacheMem_2_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2415 = 4'hf == io_writeMask ? _GEN_1903 : CacheMem_2_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2416 = 4'hf == io_writeMask ? _GEN_1904 : CacheMem_2_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2417 = 4'hf == io_writeMask ? _GEN_1905 : CacheMem_2_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2418 = 4'hf == io_writeMask ? _GEN_1906 : CacheMem_2_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2419 = 4'hf == io_writeMask ? _GEN_1907 : CacheMem_3_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2420 = 4'hf == io_writeMask ? _GEN_1908 : CacheMem_3_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2421 = 4'hf == io_writeMask ? _GEN_1909 : CacheMem_3_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2422 = 4'hf == io_writeMask ? _GEN_1910 : CacheMem_3_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2423 = 4'hf == io_writeMask ? _GEN_1911 : CacheMem_3_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2424 = 4'hf == io_writeMask ? _GEN_1912 : CacheMem_3_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2425 = 4'hf == io_writeMask ? _GEN_1913 : CacheMem_3_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2426 = 4'hf == io_writeMask ? _GEN_1914 : CacheMem_3_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2427 = 4'hf == io_writeMask ? _GEN_1915 : CacheMem_3_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2428 = 4'hf == io_writeMask ? _GEN_1916 : CacheMem_3_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2429 = 4'hf == io_writeMask ? _GEN_1917 : CacheMem_3_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2430 = 4'hf == io_writeMask ? _GEN_1918 : CacheMem_3_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2431 = 4'hf == io_writeMask ? _GEN_1919 : CacheMem_3_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2432 = 4'hf == io_writeMask ? _GEN_1920 : CacheMem_3_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2433 = 4'hf == io_writeMask ? _GEN_1921 : CacheMem_3_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2434 = 4'hf == io_writeMask ? _GEN_1922 : CacheMem_3_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2435 = 4'hf == io_writeMask ? _GEN_1923 : CacheMem_3_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2436 = 4'hf == io_writeMask ? _GEN_1924 : CacheMem_3_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2437 = 4'hf == io_writeMask ? _GEN_1925 : CacheMem_3_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2438 = 4'hf == io_writeMask ? _GEN_1926 : CacheMem_3_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2439 = 4'hf == io_writeMask ? _GEN_1927 : CacheMem_3_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2440 = 4'hf == io_writeMask ? _GEN_1928 : CacheMem_3_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2441 = 4'hf == io_writeMask ? _GEN_1929 : CacheMem_3_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2442 = 4'hf == io_writeMask ? _GEN_1930 : CacheMem_3_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2443 = 4'hf == io_writeMask ? _GEN_1931 : CacheMem_3_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2444 = 4'hf == io_writeMask ? _GEN_1932 : CacheMem_3_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2445 = 4'hf == io_writeMask ? _GEN_1933 : CacheMem_3_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2446 = 4'hf == io_writeMask ? _GEN_1934 : CacheMem_3_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2447 = 4'hf == io_writeMask ? _GEN_1935 : CacheMem_3_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2448 = 4'hf == io_writeMask ? _GEN_1936 : CacheMem_3_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2449 = 4'hf == io_writeMask ? _GEN_1937 : CacheMem_3_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2450 = 4'hf == io_writeMask ? _GEN_1938 : CacheMem_3_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2451 = 4'hf == io_writeMask ? _GEN_1939 : CacheMem_3_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2452 = 4'hf == io_writeMask ? _GEN_1940 : CacheMem_3_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2453 = 4'hf == io_writeMask ? _GEN_1941 : CacheMem_3_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2454 = 4'hf == io_writeMask ? _GEN_1942 : CacheMem_3_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2455 = 4'hf == io_writeMask ? _GEN_1943 : CacheMem_3_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2456 = 4'hf == io_writeMask ? _GEN_1944 : CacheMem_3_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2457 = 4'hf == io_writeMask ? _GEN_1945 : CacheMem_3_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2458 = 4'hf == io_writeMask ? _GEN_1946 : CacheMem_3_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2459 = 4'hf == io_writeMask ? _GEN_1947 : CacheMem_3_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2460 = 4'hf == io_writeMask ? _GEN_1948 : CacheMem_3_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2461 = 4'hf == io_writeMask ? _GEN_1949 : CacheMem_3_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2462 = 4'hf == io_writeMask ? _GEN_1950 : CacheMem_3_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2463 = 4'hf == io_writeMask ? _GEN_1951 : CacheMem_3_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2464 = 4'hf == io_writeMask ? _GEN_1952 : CacheMem_3_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2465 = 4'hf == io_writeMask ? _GEN_1953 : CacheMem_3_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2466 = 4'hf == io_writeMask ? _GEN_1954 : CacheMem_3_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2467 = 4'hf == io_writeMask ? _GEN_1955 : CacheMem_3_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2468 = 4'hf == io_writeMask ? _GEN_1956 : CacheMem_3_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2469 = 4'hf == io_writeMask ? _GEN_1957 : CacheMem_3_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2470 = 4'hf == io_writeMask ? _GEN_1958 : CacheMem_3_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2471 = 4'hf == io_writeMask ? _GEN_1959 : CacheMem_3_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2472 = 4'hf == io_writeMask ? _GEN_1960 : CacheMem_3_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2473 = 4'hf == io_writeMask ? _GEN_1961 : CacheMem_3_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2474 = 4'hf == io_writeMask ? _GEN_1962 : CacheMem_3_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2475 = 4'hf == io_writeMask ? _GEN_1963 : CacheMem_3_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2476 = 4'hf == io_writeMask ? _GEN_1964 : CacheMem_3_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2477 = 4'hf == io_writeMask ? _GEN_1965 : CacheMem_3_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2478 = 4'hf == io_writeMask ? _GEN_1966 : CacheMem_3_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2479 = 4'hf == io_writeMask ? _GEN_1967 : CacheMem_3_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2480 = 4'hf == io_writeMask ? _GEN_1968 : CacheMem_3_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2481 = 4'hf == io_writeMask ? _GEN_1969 : CacheMem_3_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2482 = 4'hf == io_writeMask ? _GEN_1970 : CacheMem_3_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2483 = 4'hf == io_writeMask ? _GEN_1971 : CacheMem_4_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2484 = 4'hf == io_writeMask ? _GEN_1972 : CacheMem_4_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2485 = 4'hf == io_writeMask ? _GEN_1973 : CacheMem_4_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2486 = 4'hf == io_writeMask ? _GEN_1974 : CacheMem_4_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2487 = 4'hf == io_writeMask ? _GEN_1975 : CacheMem_4_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2488 = 4'hf == io_writeMask ? _GEN_1976 : CacheMem_4_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2489 = 4'hf == io_writeMask ? _GEN_1977 : CacheMem_4_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2490 = 4'hf == io_writeMask ? _GEN_1978 : CacheMem_4_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2491 = 4'hf == io_writeMask ? _GEN_1979 : CacheMem_4_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2492 = 4'hf == io_writeMask ? _GEN_1980 : CacheMem_4_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2493 = 4'hf == io_writeMask ? _GEN_1981 : CacheMem_4_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2494 = 4'hf == io_writeMask ? _GEN_1982 : CacheMem_4_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2495 = 4'hf == io_writeMask ? _GEN_1983 : CacheMem_4_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2496 = 4'hf == io_writeMask ? _GEN_1984 : CacheMem_4_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2497 = 4'hf == io_writeMask ? _GEN_1985 : CacheMem_4_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2498 = 4'hf == io_writeMask ? _GEN_1986 : CacheMem_4_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2499 = 4'hf == io_writeMask ? _GEN_1987 : CacheMem_4_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2500 = 4'hf == io_writeMask ? _GEN_1988 : CacheMem_4_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2501 = 4'hf == io_writeMask ? _GEN_1989 : CacheMem_4_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2502 = 4'hf == io_writeMask ? _GEN_1990 : CacheMem_4_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2503 = 4'hf == io_writeMask ? _GEN_1991 : CacheMem_4_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2504 = 4'hf == io_writeMask ? _GEN_1992 : CacheMem_4_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2505 = 4'hf == io_writeMask ? _GEN_1993 : CacheMem_4_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2506 = 4'hf == io_writeMask ? _GEN_1994 : CacheMem_4_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2507 = 4'hf == io_writeMask ? _GEN_1995 : CacheMem_4_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2508 = 4'hf == io_writeMask ? _GEN_1996 : CacheMem_4_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2509 = 4'hf == io_writeMask ? _GEN_1997 : CacheMem_4_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2510 = 4'hf == io_writeMask ? _GEN_1998 : CacheMem_4_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2511 = 4'hf == io_writeMask ? _GEN_1999 : CacheMem_4_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2512 = 4'hf == io_writeMask ? _GEN_2000 : CacheMem_4_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2513 = 4'hf == io_writeMask ? _GEN_2001 : CacheMem_4_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2514 = 4'hf == io_writeMask ? _GEN_2002 : CacheMem_4_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2515 = 4'hf == io_writeMask ? _GEN_2003 : CacheMem_4_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2516 = 4'hf == io_writeMask ? _GEN_2004 : CacheMem_4_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2517 = 4'hf == io_writeMask ? _GEN_2005 : CacheMem_4_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2518 = 4'hf == io_writeMask ? _GEN_2006 : CacheMem_4_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2519 = 4'hf == io_writeMask ? _GEN_2007 : CacheMem_4_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2520 = 4'hf == io_writeMask ? _GEN_2008 : CacheMem_4_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2521 = 4'hf == io_writeMask ? _GEN_2009 : CacheMem_4_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2522 = 4'hf == io_writeMask ? _GEN_2010 : CacheMem_4_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2523 = 4'hf == io_writeMask ? _GEN_2011 : CacheMem_4_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2524 = 4'hf == io_writeMask ? _GEN_2012 : CacheMem_4_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2525 = 4'hf == io_writeMask ? _GEN_2013 : CacheMem_4_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2526 = 4'hf == io_writeMask ? _GEN_2014 : CacheMem_4_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2527 = 4'hf == io_writeMask ? _GEN_2015 : CacheMem_4_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2528 = 4'hf == io_writeMask ? _GEN_2016 : CacheMem_4_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2529 = 4'hf == io_writeMask ? _GEN_2017 : CacheMem_4_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2530 = 4'hf == io_writeMask ? _GEN_2018 : CacheMem_4_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2531 = 4'hf == io_writeMask ? _GEN_2019 : CacheMem_4_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2532 = 4'hf == io_writeMask ? _GEN_2020 : CacheMem_4_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2533 = 4'hf == io_writeMask ? _GEN_2021 : CacheMem_4_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2534 = 4'hf == io_writeMask ? _GEN_2022 : CacheMem_4_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2535 = 4'hf == io_writeMask ? _GEN_2023 : CacheMem_4_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2536 = 4'hf == io_writeMask ? _GEN_2024 : CacheMem_4_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2537 = 4'hf == io_writeMask ? _GEN_2025 : CacheMem_4_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2538 = 4'hf == io_writeMask ? _GEN_2026 : CacheMem_4_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2539 = 4'hf == io_writeMask ? _GEN_2027 : CacheMem_4_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2540 = 4'hf == io_writeMask ? _GEN_2028 : CacheMem_4_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2541 = 4'hf == io_writeMask ? _GEN_2029 : CacheMem_4_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2542 = 4'hf == io_writeMask ? _GEN_2030 : CacheMem_4_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2543 = 4'hf == io_writeMask ? _GEN_2031 : CacheMem_4_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2544 = 4'hf == io_writeMask ? _GEN_2032 : CacheMem_4_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2545 = 4'hf == io_writeMask ? _GEN_2033 : CacheMem_4_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2546 = 4'hf == io_writeMask ? _GEN_2034 : CacheMem_4_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2547 = 4'hf == io_writeMask ? _GEN_2035 : CacheMem_5_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2548 = 4'hf == io_writeMask ? _GEN_2036 : CacheMem_5_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2549 = 4'hf == io_writeMask ? _GEN_2037 : CacheMem_5_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2550 = 4'hf == io_writeMask ? _GEN_2038 : CacheMem_5_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2551 = 4'hf == io_writeMask ? _GEN_2039 : CacheMem_5_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2552 = 4'hf == io_writeMask ? _GEN_2040 : CacheMem_5_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2553 = 4'hf == io_writeMask ? _GEN_2041 : CacheMem_5_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2554 = 4'hf == io_writeMask ? _GEN_2042 : CacheMem_5_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2555 = 4'hf == io_writeMask ? _GEN_2043 : CacheMem_5_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2556 = 4'hf == io_writeMask ? _GEN_2044 : CacheMem_5_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2557 = 4'hf == io_writeMask ? _GEN_2045 : CacheMem_5_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2558 = 4'hf == io_writeMask ? _GEN_2046 : CacheMem_5_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2559 = 4'hf == io_writeMask ? _GEN_2047 : CacheMem_5_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2560 = 4'hf == io_writeMask ? _GEN_2048 : CacheMem_5_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2561 = 4'hf == io_writeMask ? _GEN_2049 : CacheMem_5_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2562 = 4'hf == io_writeMask ? _GEN_2050 : CacheMem_5_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2563 = 4'hf == io_writeMask ? _GEN_2051 : CacheMem_5_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2564 = 4'hf == io_writeMask ? _GEN_2052 : CacheMem_5_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2565 = 4'hf == io_writeMask ? _GEN_2053 : CacheMem_5_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2566 = 4'hf == io_writeMask ? _GEN_2054 : CacheMem_5_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2567 = 4'hf == io_writeMask ? _GEN_2055 : CacheMem_5_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2568 = 4'hf == io_writeMask ? _GEN_2056 : CacheMem_5_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2569 = 4'hf == io_writeMask ? _GEN_2057 : CacheMem_5_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2570 = 4'hf == io_writeMask ? _GEN_2058 : CacheMem_5_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2571 = 4'hf == io_writeMask ? _GEN_2059 : CacheMem_5_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2572 = 4'hf == io_writeMask ? _GEN_2060 : CacheMem_5_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2573 = 4'hf == io_writeMask ? _GEN_2061 : CacheMem_5_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2574 = 4'hf == io_writeMask ? _GEN_2062 : CacheMem_5_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2575 = 4'hf == io_writeMask ? _GEN_2063 : CacheMem_5_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2576 = 4'hf == io_writeMask ? _GEN_2064 : CacheMem_5_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2577 = 4'hf == io_writeMask ? _GEN_2065 : CacheMem_5_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2578 = 4'hf == io_writeMask ? _GEN_2066 : CacheMem_5_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2579 = 4'hf == io_writeMask ? _GEN_2067 : CacheMem_5_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2580 = 4'hf == io_writeMask ? _GEN_2068 : CacheMem_5_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2581 = 4'hf == io_writeMask ? _GEN_2069 : CacheMem_5_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2582 = 4'hf == io_writeMask ? _GEN_2070 : CacheMem_5_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2583 = 4'hf == io_writeMask ? _GEN_2071 : CacheMem_5_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2584 = 4'hf == io_writeMask ? _GEN_2072 : CacheMem_5_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2585 = 4'hf == io_writeMask ? _GEN_2073 : CacheMem_5_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2586 = 4'hf == io_writeMask ? _GEN_2074 : CacheMem_5_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2587 = 4'hf == io_writeMask ? _GEN_2075 : CacheMem_5_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2588 = 4'hf == io_writeMask ? _GEN_2076 : CacheMem_5_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2589 = 4'hf == io_writeMask ? _GEN_2077 : CacheMem_5_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2590 = 4'hf == io_writeMask ? _GEN_2078 : CacheMem_5_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2591 = 4'hf == io_writeMask ? _GEN_2079 : CacheMem_5_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2592 = 4'hf == io_writeMask ? _GEN_2080 : CacheMem_5_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2593 = 4'hf == io_writeMask ? _GEN_2081 : CacheMem_5_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2594 = 4'hf == io_writeMask ? _GEN_2082 : CacheMem_5_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2595 = 4'hf == io_writeMask ? _GEN_2083 : CacheMem_5_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2596 = 4'hf == io_writeMask ? _GEN_2084 : CacheMem_5_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2597 = 4'hf == io_writeMask ? _GEN_2085 : CacheMem_5_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2598 = 4'hf == io_writeMask ? _GEN_2086 : CacheMem_5_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2599 = 4'hf == io_writeMask ? _GEN_2087 : CacheMem_5_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2600 = 4'hf == io_writeMask ? _GEN_2088 : CacheMem_5_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2601 = 4'hf == io_writeMask ? _GEN_2089 : CacheMem_5_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2602 = 4'hf == io_writeMask ? _GEN_2090 : CacheMem_5_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2603 = 4'hf == io_writeMask ? _GEN_2091 : CacheMem_5_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2604 = 4'hf == io_writeMask ? _GEN_2092 : CacheMem_5_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2605 = 4'hf == io_writeMask ? _GEN_2093 : CacheMem_5_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2606 = 4'hf == io_writeMask ? _GEN_2094 : CacheMem_5_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2607 = 4'hf == io_writeMask ? _GEN_2095 : CacheMem_5_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2608 = 4'hf == io_writeMask ? _GEN_2096 : CacheMem_5_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2609 = 4'hf == io_writeMask ? _GEN_2097 : CacheMem_5_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2610 = 4'hf == io_writeMask ? _GEN_2098 : CacheMem_5_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2611 = 4'hf == io_writeMask ? _GEN_2099 : CacheMem_6_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2612 = 4'hf == io_writeMask ? _GEN_2100 : CacheMem_6_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2613 = 4'hf == io_writeMask ? _GEN_2101 : CacheMem_6_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2614 = 4'hf == io_writeMask ? _GEN_2102 : CacheMem_6_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2615 = 4'hf == io_writeMask ? _GEN_2103 : CacheMem_6_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2616 = 4'hf == io_writeMask ? _GEN_2104 : CacheMem_6_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2617 = 4'hf == io_writeMask ? _GEN_2105 : CacheMem_6_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2618 = 4'hf == io_writeMask ? _GEN_2106 : CacheMem_6_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2619 = 4'hf == io_writeMask ? _GEN_2107 : CacheMem_6_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2620 = 4'hf == io_writeMask ? _GEN_2108 : CacheMem_6_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2621 = 4'hf == io_writeMask ? _GEN_2109 : CacheMem_6_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2622 = 4'hf == io_writeMask ? _GEN_2110 : CacheMem_6_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2623 = 4'hf == io_writeMask ? _GEN_2111 : CacheMem_6_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2624 = 4'hf == io_writeMask ? _GEN_2112 : CacheMem_6_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2625 = 4'hf == io_writeMask ? _GEN_2113 : CacheMem_6_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2626 = 4'hf == io_writeMask ? _GEN_2114 : CacheMem_6_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2627 = 4'hf == io_writeMask ? _GEN_2115 : CacheMem_6_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2628 = 4'hf == io_writeMask ? _GEN_2116 : CacheMem_6_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2629 = 4'hf == io_writeMask ? _GEN_2117 : CacheMem_6_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2630 = 4'hf == io_writeMask ? _GEN_2118 : CacheMem_6_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2631 = 4'hf == io_writeMask ? _GEN_2119 : CacheMem_6_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2632 = 4'hf == io_writeMask ? _GEN_2120 : CacheMem_6_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2633 = 4'hf == io_writeMask ? _GEN_2121 : CacheMem_6_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2634 = 4'hf == io_writeMask ? _GEN_2122 : CacheMem_6_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2635 = 4'hf == io_writeMask ? _GEN_2123 : CacheMem_6_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2636 = 4'hf == io_writeMask ? _GEN_2124 : CacheMem_6_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2637 = 4'hf == io_writeMask ? _GEN_2125 : CacheMem_6_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2638 = 4'hf == io_writeMask ? _GEN_2126 : CacheMem_6_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2639 = 4'hf == io_writeMask ? _GEN_2127 : CacheMem_6_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2640 = 4'hf == io_writeMask ? _GEN_2128 : CacheMem_6_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2641 = 4'hf == io_writeMask ? _GEN_2129 : CacheMem_6_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2642 = 4'hf == io_writeMask ? _GEN_2130 : CacheMem_6_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2643 = 4'hf == io_writeMask ? _GEN_2131 : CacheMem_6_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2644 = 4'hf == io_writeMask ? _GEN_2132 : CacheMem_6_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2645 = 4'hf == io_writeMask ? _GEN_2133 : CacheMem_6_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2646 = 4'hf == io_writeMask ? _GEN_2134 : CacheMem_6_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2647 = 4'hf == io_writeMask ? _GEN_2135 : CacheMem_6_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2648 = 4'hf == io_writeMask ? _GEN_2136 : CacheMem_6_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2649 = 4'hf == io_writeMask ? _GEN_2137 : CacheMem_6_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2650 = 4'hf == io_writeMask ? _GEN_2138 : CacheMem_6_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2651 = 4'hf == io_writeMask ? _GEN_2139 : CacheMem_6_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2652 = 4'hf == io_writeMask ? _GEN_2140 : CacheMem_6_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2653 = 4'hf == io_writeMask ? _GEN_2141 : CacheMem_6_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2654 = 4'hf == io_writeMask ? _GEN_2142 : CacheMem_6_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2655 = 4'hf == io_writeMask ? _GEN_2143 : CacheMem_6_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2656 = 4'hf == io_writeMask ? _GEN_2144 : CacheMem_6_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2657 = 4'hf == io_writeMask ? _GEN_2145 : CacheMem_6_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2658 = 4'hf == io_writeMask ? _GEN_2146 : CacheMem_6_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2659 = 4'hf == io_writeMask ? _GEN_2147 : CacheMem_6_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2660 = 4'hf == io_writeMask ? _GEN_2148 : CacheMem_6_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2661 = 4'hf == io_writeMask ? _GEN_2149 : CacheMem_6_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2662 = 4'hf == io_writeMask ? _GEN_2150 : CacheMem_6_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2663 = 4'hf == io_writeMask ? _GEN_2151 : CacheMem_6_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2664 = 4'hf == io_writeMask ? _GEN_2152 : CacheMem_6_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2665 = 4'hf == io_writeMask ? _GEN_2153 : CacheMem_6_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2666 = 4'hf == io_writeMask ? _GEN_2154 : CacheMem_6_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2667 = 4'hf == io_writeMask ? _GEN_2155 : CacheMem_6_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2668 = 4'hf == io_writeMask ? _GEN_2156 : CacheMem_6_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2669 = 4'hf == io_writeMask ? _GEN_2157 : CacheMem_6_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2670 = 4'hf == io_writeMask ? _GEN_2158 : CacheMem_6_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2671 = 4'hf == io_writeMask ? _GEN_2159 : CacheMem_6_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2672 = 4'hf == io_writeMask ? _GEN_2160 : CacheMem_6_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2673 = 4'hf == io_writeMask ? _GEN_2161 : CacheMem_6_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2674 = 4'hf == io_writeMask ? _GEN_2162 : CacheMem_6_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2675 = 4'hf == io_writeMask ? _GEN_2163 : CacheMem_7_0_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2676 = 4'hf == io_writeMask ? _GEN_2164 : CacheMem_7_0_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2677 = 4'hf == io_writeMask ? _GEN_2165 : CacheMem_7_0_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2678 = 4'hf == io_writeMask ? _GEN_2166 : CacheMem_7_0_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2679 = 4'hf == io_writeMask ? _GEN_2167 : CacheMem_7_0_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2680 = 4'hf == io_writeMask ? _GEN_2168 : CacheMem_7_0_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2681 = 4'hf == io_writeMask ? _GEN_2169 : CacheMem_7_0_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2682 = 4'hf == io_writeMask ? _GEN_2170 : CacheMem_7_0_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2683 = 4'hf == io_writeMask ? _GEN_2171 : CacheMem_7_1_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2684 = 4'hf == io_writeMask ? _GEN_2172 : CacheMem_7_1_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2685 = 4'hf == io_writeMask ? _GEN_2173 : CacheMem_7_1_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2686 = 4'hf == io_writeMask ? _GEN_2174 : CacheMem_7_1_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2687 = 4'hf == io_writeMask ? _GEN_2175 : CacheMem_7_1_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2688 = 4'hf == io_writeMask ? _GEN_2176 : CacheMem_7_1_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2689 = 4'hf == io_writeMask ? _GEN_2177 : CacheMem_7_1_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2690 = 4'hf == io_writeMask ? _GEN_2178 : CacheMem_7_1_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2691 = 4'hf == io_writeMask ? _GEN_2179 : CacheMem_7_2_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2692 = 4'hf == io_writeMask ? _GEN_2180 : CacheMem_7_2_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2693 = 4'hf == io_writeMask ? _GEN_2181 : CacheMem_7_2_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2694 = 4'hf == io_writeMask ? _GEN_2182 : CacheMem_7_2_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2695 = 4'hf == io_writeMask ? _GEN_2183 : CacheMem_7_2_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2696 = 4'hf == io_writeMask ? _GEN_2184 : CacheMem_7_2_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2697 = 4'hf == io_writeMask ? _GEN_2185 : CacheMem_7_2_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2698 = 4'hf == io_writeMask ? _GEN_2186 : CacheMem_7_2_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2699 = 4'hf == io_writeMask ? _GEN_2187 : CacheMem_7_3_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2700 = 4'hf == io_writeMask ? _GEN_2188 : CacheMem_7_3_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2701 = 4'hf == io_writeMask ? _GEN_2189 : CacheMem_7_3_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2702 = 4'hf == io_writeMask ? _GEN_2190 : CacheMem_7_3_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2703 = 4'hf == io_writeMask ? _GEN_2191 : CacheMem_7_3_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2704 = 4'hf == io_writeMask ? _GEN_2192 : CacheMem_7_3_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2705 = 4'hf == io_writeMask ? _GEN_2193 : CacheMem_7_3_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2706 = 4'hf == io_writeMask ? _GEN_2194 : CacheMem_7_3_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2707 = 4'hf == io_writeMask ? _GEN_2195 : CacheMem_7_4_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2708 = 4'hf == io_writeMask ? _GEN_2196 : CacheMem_7_4_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2709 = 4'hf == io_writeMask ? _GEN_2197 : CacheMem_7_4_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2710 = 4'hf == io_writeMask ? _GEN_2198 : CacheMem_7_4_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2711 = 4'hf == io_writeMask ? _GEN_2199 : CacheMem_7_4_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2712 = 4'hf == io_writeMask ? _GEN_2200 : CacheMem_7_4_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2713 = 4'hf == io_writeMask ? _GEN_2201 : CacheMem_7_4_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2714 = 4'hf == io_writeMask ? _GEN_2202 : CacheMem_7_4_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2715 = 4'hf == io_writeMask ? _GEN_2203 : CacheMem_7_5_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2716 = 4'hf == io_writeMask ? _GEN_2204 : CacheMem_7_5_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2717 = 4'hf == io_writeMask ? _GEN_2205 : CacheMem_7_5_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2718 = 4'hf == io_writeMask ? _GEN_2206 : CacheMem_7_5_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2719 = 4'hf == io_writeMask ? _GEN_2207 : CacheMem_7_5_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2720 = 4'hf == io_writeMask ? _GEN_2208 : CacheMem_7_5_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2721 = 4'hf == io_writeMask ? _GEN_2209 : CacheMem_7_5_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2722 = 4'hf == io_writeMask ? _GEN_2210 : CacheMem_7_5_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2723 = 4'hf == io_writeMask ? _GEN_2211 : CacheMem_7_6_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2724 = 4'hf == io_writeMask ? _GEN_2212 : CacheMem_7_6_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2725 = 4'hf == io_writeMask ? _GEN_2213 : CacheMem_7_6_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2726 = 4'hf == io_writeMask ? _GEN_2214 : CacheMem_7_6_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2727 = 4'hf == io_writeMask ? _GEN_2215 : CacheMem_7_6_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2728 = 4'hf == io_writeMask ? _GEN_2216 : CacheMem_7_6_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2729 = 4'hf == io_writeMask ? _GEN_2217 : CacheMem_7_6_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2730 = 4'hf == io_writeMask ? _GEN_2218 : CacheMem_7_6_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2731 = 4'hf == io_writeMask ? _GEN_2219 : CacheMem_7_7_0; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2732 = 4'hf == io_writeMask ? _GEN_2220 : CacheMem_7_7_1; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2733 = 4'hf == io_writeMask ? _GEN_2221 : CacheMem_7_7_2; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2734 = 4'hf == io_writeMask ? _GEN_2222 : CacheMem_7_7_3; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2735 = 4'hf == io_writeMask ? _GEN_2223 : CacheMem_7_7_4; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2736 = 4'hf == io_writeMask ? _GEN_2224 : CacheMem_7_7_5; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2737 = 4'hf == io_writeMask ? _GEN_2225 : CacheMem_7_7_6; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2738 = 4'hf == io_writeMask ? _GEN_2226 : CacheMem_7_7_7; // @[Cache.scala 133:31 53:25]
  wire [31:0] _GEN_2739 = 4'h3 == io_writeMask ? _GEN_1203 : _GEN_2227; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2740 = 4'h3 == io_writeMask ? _GEN_1204 : _GEN_2228; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2741 = 4'h3 == io_writeMask ? _GEN_1205 : _GEN_2229; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2742 = 4'h3 == io_writeMask ? _GEN_1206 : _GEN_2230; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2743 = 4'h3 == io_writeMask ? _GEN_1207 : _GEN_2231; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2744 = 4'h3 == io_writeMask ? _GEN_1208 : _GEN_2232; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2745 = 4'h3 == io_writeMask ? _GEN_1209 : _GEN_2233; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2746 = 4'h3 == io_writeMask ? _GEN_1210 : _GEN_2234; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2747 = 4'h3 == io_writeMask ? _GEN_1211 : _GEN_2235; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2748 = 4'h3 == io_writeMask ? _GEN_1212 : _GEN_2236; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2749 = 4'h3 == io_writeMask ? _GEN_1213 : _GEN_2237; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2750 = 4'h3 == io_writeMask ? _GEN_1214 : _GEN_2238; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2751 = 4'h3 == io_writeMask ? _GEN_1215 : _GEN_2239; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2752 = 4'h3 == io_writeMask ? _GEN_1216 : _GEN_2240; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2753 = 4'h3 == io_writeMask ? _GEN_1217 : _GEN_2241; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2754 = 4'h3 == io_writeMask ? _GEN_1218 : _GEN_2242; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2755 = 4'h3 == io_writeMask ? _GEN_1219 : _GEN_2243; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2756 = 4'h3 == io_writeMask ? _GEN_1220 : _GEN_2244; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2757 = 4'h3 == io_writeMask ? _GEN_1221 : _GEN_2245; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2758 = 4'h3 == io_writeMask ? _GEN_1222 : _GEN_2246; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2759 = 4'h3 == io_writeMask ? _GEN_1223 : _GEN_2247; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2760 = 4'h3 == io_writeMask ? _GEN_1224 : _GEN_2248; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2761 = 4'h3 == io_writeMask ? _GEN_1225 : _GEN_2249; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2762 = 4'h3 == io_writeMask ? _GEN_1226 : _GEN_2250; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2763 = 4'h3 == io_writeMask ? _GEN_1227 : _GEN_2251; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2764 = 4'h3 == io_writeMask ? _GEN_1228 : _GEN_2252; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2765 = 4'h3 == io_writeMask ? _GEN_1229 : _GEN_2253; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2766 = 4'h3 == io_writeMask ? _GEN_1230 : _GEN_2254; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2767 = 4'h3 == io_writeMask ? _GEN_1231 : _GEN_2255; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2768 = 4'h3 == io_writeMask ? _GEN_1232 : _GEN_2256; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2769 = 4'h3 == io_writeMask ? _GEN_1233 : _GEN_2257; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2770 = 4'h3 == io_writeMask ? _GEN_1234 : _GEN_2258; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2771 = 4'h3 == io_writeMask ? _GEN_1235 : _GEN_2259; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2772 = 4'h3 == io_writeMask ? _GEN_1236 : _GEN_2260; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2773 = 4'h3 == io_writeMask ? _GEN_1237 : _GEN_2261; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2774 = 4'h3 == io_writeMask ? _GEN_1238 : _GEN_2262; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2775 = 4'h3 == io_writeMask ? _GEN_1239 : _GEN_2263; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2776 = 4'h3 == io_writeMask ? _GEN_1240 : _GEN_2264; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2777 = 4'h3 == io_writeMask ? _GEN_1241 : _GEN_2265; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2778 = 4'h3 == io_writeMask ? _GEN_1242 : _GEN_2266; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2779 = 4'h3 == io_writeMask ? _GEN_1243 : _GEN_2267; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2780 = 4'h3 == io_writeMask ? _GEN_1244 : _GEN_2268; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2781 = 4'h3 == io_writeMask ? _GEN_1245 : _GEN_2269; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2782 = 4'h3 == io_writeMask ? _GEN_1246 : _GEN_2270; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2783 = 4'h3 == io_writeMask ? _GEN_1247 : _GEN_2271; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2784 = 4'h3 == io_writeMask ? _GEN_1248 : _GEN_2272; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2785 = 4'h3 == io_writeMask ? _GEN_1249 : _GEN_2273; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2786 = 4'h3 == io_writeMask ? _GEN_1250 : _GEN_2274; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2787 = 4'h3 == io_writeMask ? _GEN_1251 : _GEN_2275; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2788 = 4'h3 == io_writeMask ? _GEN_1252 : _GEN_2276; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2789 = 4'h3 == io_writeMask ? _GEN_1253 : _GEN_2277; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2790 = 4'h3 == io_writeMask ? _GEN_1254 : _GEN_2278; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2791 = 4'h3 == io_writeMask ? _GEN_1255 : _GEN_2279; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2792 = 4'h3 == io_writeMask ? _GEN_1256 : _GEN_2280; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2793 = 4'h3 == io_writeMask ? _GEN_1257 : _GEN_2281; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2794 = 4'h3 == io_writeMask ? _GEN_1258 : _GEN_2282; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2795 = 4'h3 == io_writeMask ? _GEN_1259 : _GEN_2283; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2796 = 4'h3 == io_writeMask ? _GEN_1260 : _GEN_2284; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2797 = 4'h3 == io_writeMask ? _GEN_1261 : _GEN_2285; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2798 = 4'h3 == io_writeMask ? _GEN_1262 : _GEN_2286; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2799 = 4'h3 == io_writeMask ? _GEN_1263 : _GEN_2287; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2800 = 4'h3 == io_writeMask ? _GEN_1264 : _GEN_2288; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2801 = 4'h3 == io_writeMask ? _GEN_1265 : _GEN_2289; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2802 = 4'h3 == io_writeMask ? _GEN_1266 : _GEN_2290; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2803 = 4'h3 == io_writeMask ? _GEN_1267 : _GEN_2291; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2804 = 4'h3 == io_writeMask ? _GEN_1268 : _GEN_2292; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2805 = 4'h3 == io_writeMask ? _GEN_1269 : _GEN_2293; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2806 = 4'h3 == io_writeMask ? _GEN_1270 : _GEN_2294; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2807 = 4'h3 == io_writeMask ? _GEN_1271 : _GEN_2295; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2808 = 4'h3 == io_writeMask ? _GEN_1272 : _GEN_2296; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2809 = 4'h3 == io_writeMask ? _GEN_1273 : _GEN_2297; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2810 = 4'h3 == io_writeMask ? _GEN_1274 : _GEN_2298; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2811 = 4'h3 == io_writeMask ? _GEN_1275 : _GEN_2299; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2812 = 4'h3 == io_writeMask ? _GEN_1276 : _GEN_2300; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2813 = 4'h3 == io_writeMask ? _GEN_1277 : _GEN_2301; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2814 = 4'h3 == io_writeMask ? _GEN_1278 : _GEN_2302; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2815 = 4'h3 == io_writeMask ? _GEN_1279 : _GEN_2303; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2816 = 4'h3 == io_writeMask ? _GEN_1280 : _GEN_2304; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2817 = 4'h3 == io_writeMask ? _GEN_1281 : _GEN_2305; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2818 = 4'h3 == io_writeMask ? _GEN_1282 : _GEN_2306; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2819 = 4'h3 == io_writeMask ? _GEN_1283 : _GEN_2307; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2820 = 4'h3 == io_writeMask ? _GEN_1284 : _GEN_2308; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2821 = 4'h3 == io_writeMask ? _GEN_1285 : _GEN_2309; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2822 = 4'h3 == io_writeMask ? _GEN_1286 : _GEN_2310; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2823 = 4'h3 == io_writeMask ? _GEN_1287 : _GEN_2311; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2824 = 4'h3 == io_writeMask ? _GEN_1288 : _GEN_2312; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2825 = 4'h3 == io_writeMask ? _GEN_1289 : _GEN_2313; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2826 = 4'h3 == io_writeMask ? _GEN_1290 : _GEN_2314; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2827 = 4'h3 == io_writeMask ? _GEN_1291 : _GEN_2315; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2828 = 4'h3 == io_writeMask ? _GEN_1292 : _GEN_2316; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2829 = 4'h3 == io_writeMask ? _GEN_1293 : _GEN_2317; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2830 = 4'h3 == io_writeMask ? _GEN_1294 : _GEN_2318; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2831 = 4'h3 == io_writeMask ? _GEN_1295 : _GEN_2319; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2832 = 4'h3 == io_writeMask ? _GEN_1296 : _GEN_2320; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2833 = 4'h3 == io_writeMask ? _GEN_1297 : _GEN_2321; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2834 = 4'h3 == io_writeMask ? _GEN_1298 : _GEN_2322; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2835 = 4'h3 == io_writeMask ? _GEN_1299 : _GEN_2323; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2836 = 4'h3 == io_writeMask ? _GEN_1300 : _GEN_2324; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2837 = 4'h3 == io_writeMask ? _GEN_1301 : _GEN_2325; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2838 = 4'h3 == io_writeMask ? _GEN_1302 : _GEN_2326; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2839 = 4'h3 == io_writeMask ? _GEN_1303 : _GEN_2327; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2840 = 4'h3 == io_writeMask ? _GEN_1304 : _GEN_2328; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2841 = 4'h3 == io_writeMask ? _GEN_1305 : _GEN_2329; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2842 = 4'h3 == io_writeMask ? _GEN_1306 : _GEN_2330; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2843 = 4'h3 == io_writeMask ? _GEN_1307 : _GEN_2331; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2844 = 4'h3 == io_writeMask ? _GEN_1308 : _GEN_2332; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2845 = 4'h3 == io_writeMask ? _GEN_1309 : _GEN_2333; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2846 = 4'h3 == io_writeMask ? _GEN_1310 : _GEN_2334; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2847 = 4'h3 == io_writeMask ? _GEN_1311 : _GEN_2335; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2848 = 4'h3 == io_writeMask ? _GEN_1312 : _GEN_2336; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2849 = 4'h3 == io_writeMask ? _GEN_1313 : _GEN_2337; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2850 = 4'h3 == io_writeMask ? _GEN_1314 : _GEN_2338; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2851 = 4'h3 == io_writeMask ? _GEN_1315 : _GEN_2339; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2852 = 4'h3 == io_writeMask ? _GEN_1316 : _GEN_2340; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2853 = 4'h3 == io_writeMask ? _GEN_1317 : _GEN_2341; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2854 = 4'h3 == io_writeMask ? _GEN_1318 : _GEN_2342; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2855 = 4'h3 == io_writeMask ? _GEN_1319 : _GEN_2343; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2856 = 4'h3 == io_writeMask ? _GEN_1320 : _GEN_2344; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2857 = 4'h3 == io_writeMask ? _GEN_1321 : _GEN_2345; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2858 = 4'h3 == io_writeMask ? _GEN_1322 : _GEN_2346; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2859 = 4'h3 == io_writeMask ? _GEN_1323 : _GEN_2347; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2860 = 4'h3 == io_writeMask ? _GEN_1324 : _GEN_2348; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2861 = 4'h3 == io_writeMask ? _GEN_1325 : _GEN_2349; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2862 = 4'h3 == io_writeMask ? _GEN_1326 : _GEN_2350; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2863 = 4'h3 == io_writeMask ? _GEN_1327 : _GEN_2351; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2864 = 4'h3 == io_writeMask ? _GEN_1328 : _GEN_2352; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2865 = 4'h3 == io_writeMask ? _GEN_1329 : _GEN_2353; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2866 = 4'h3 == io_writeMask ? _GEN_1330 : _GEN_2354; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2867 = 4'h3 == io_writeMask ? _GEN_1331 : _GEN_2355; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2868 = 4'h3 == io_writeMask ? _GEN_1332 : _GEN_2356; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2869 = 4'h3 == io_writeMask ? _GEN_1333 : _GEN_2357; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2870 = 4'h3 == io_writeMask ? _GEN_1334 : _GEN_2358; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2871 = 4'h3 == io_writeMask ? _GEN_1335 : _GEN_2359; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2872 = 4'h3 == io_writeMask ? _GEN_1336 : _GEN_2360; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2873 = 4'h3 == io_writeMask ? _GEN_1337 : _GEN_2361; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2874 = 4'h3 == io_writeMask ? _GEN_1338 : _GEN_2362; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2875 = 4'h3 == io_writeMask ? _GEN_1339 : _GEN_2363; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2876 = 4'h3 == io_writeMask ? _GEN_1340 : _GEN_2364; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2877 = 4'h3 == io_writeMask ? _GEN_1341 : _GEN_2365; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2878 = 4'h3 == io_writeMask ? _GEN_1342 : _GEN_2366; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2879 = 4'h3 == io_writeMask ? _GEN_1343 : _GEN_2367; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2880 = 4'h3 == io_writeMask ? _GEN_1344 : _GEN_2368; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2881 = 4'h3 == io_writeMask ? _GEN_1345 : _GEN_2369; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2882 = 4'h3 == io_writeMask ? _GEN_1346 : _GEN_2370; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2883 = 4'h3 == io_writeMask ? _GEN_1347 : _GEN_2371; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2884 = 4'h3 == io_writeMask ? _GEN_1348 : _GEN_2372; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2885 = 4'h3 == io_writeMask ? _GEN_1349 : _GEN_2373; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2886 = 4'h3 == io_writeMask ? _GEN_1350 : _GEN_2374; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2887 = 4'h3 == io_writeMask ? _GEN_1351 : _GEN_2375; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2888 = 4'h3 == io_writeMask ? _GEN_1352 : _GEN_2376; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2889 = 4'h3 == io_writeMask ? _GEN_1353 : _GEN_2377; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2890 = 4'h3 == io_writeMask ? _GEN_1354 : _GEN_2378; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2891 = 4'h3 == io_writeMask ? _GEN_1355 : _GEN_2379; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2892 = 4'h3 == io_writeMask ? _GEN_1356 : _GEN_2380; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2893 = 4'h3 == io_writeMask ? _GEN_1357 : _GEN_2381; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2894 = 4'h3 == io_writeMask ? _GEN_1358 : _GEN_2382; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2895 = 4'h3 == io_writeMask ? _GEN_1359 : _GEN_2383; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2896 = 4'h3 == io_writeMask ? _GEN_1360 : _GEN_2384; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2897 = 4'h3 == io_writeMask ? _GEN_1361 : _GEN_2385; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2898 = 4'h3 == io_writeMask ? _GEN_1362 : _GEN_2386; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2899 = 4'h3 == io_writeMask ? _GEN_1363 : _GEN_2387; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2900 = 4'h3 == io_writeMask ? _GEN_1364 : _GEN_2388; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2901 = 4'h3 == io_writeMask ? _GEN_1365 : _GEN_2389; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2902 = 4'h3 == io_writeMask ? _GEN_1366 : _GEN_2390; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2903 = 4'h3 == io_writeMask ? _GEN_1367 : _GEN_2391; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2904 = 4'h3 == io_writeMask ? _GEN_1368 : _GEN_2392; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2905 = 4'h3 == io_writeMask ? _GEN_1369 : _GEN_2393; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2906 = 4'h3 == io_writeMask ? _GEN_1370 : _GEN_2394; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2907 = 4'h3 == io_writeMask ? _GEN_1371 : _GEN_2395; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2908 = 4'h3 == io_writeMask ? _GEN_1372 : _GEN_2396; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2909 = 4'h3 == io_writeMask ? _GEN_1373 : _GEN_2397; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2910 = 4'h3 == io_writeMask ? _GEN_1374 : _GEN_2398; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2911 = 4'h3 == io_writeMask ? _GEN_1375 : _GEN_2399; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2912 = 4'h3 == io_writeMask ? _GEN_1376 : _GEN_2400; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2913 = 4'h3 == io_writeMask ? _GEN_1377 : _GEN_2401; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2914 = 4'h3 == io_writeMask ? _GEN_1378 : _GEN_2402; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2915 = 4'h3 == io_writeMask ? _GEN_1379 : _GEN_2403; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2916 = 4'h3 == io_writeMask ? _GEN_1380 : _GEN_2404; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2917 = 4'h3 == io_writeMask ? _GEN_1381 : _GEN_2405; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2918 = 4'h3 == io_writeMask ? _GEN_1382 : _GEN_2406; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2919 = 4'h3 == io_writeMask ? _GEN_1383 : _GEN_2407; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2920 = 4'h3 == io_writeMask ? _GEN_1384 : _GEN_2408; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2921 = 4'h3 == io_writeMask ? _GEN_1385 : _GEN_2409; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2922 = 4'h3 == io_writeMask ? _GEN_1386 : _GEN_2410; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2923 = 4'h3 == io_writeMask ? _GEN_1387 : _GEN_2411; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2924 = 4'h3 == io_writeMask ? _GEN_1388 : _GEN_2412; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2925 = 4'h3 == io_writeMask ? _GEN_1389 : _GEN_2413; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2926 = 4'h3 == io_writeMask ? _GEN_1390 : _GEN_2414; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2927 = 4'h3 == io_writeMask ? _GEN_1391 : _GEN_2415; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2928 = 4'h3 == io_writeMask ? _GEN_1392 : _GEN_2416; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2929 = 4'h3 == io_writeMask ? _GEN_1393 : _GEN_2417; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2930 = 4'h3 == io_writeMask ? _GEN_1394 : _GEN_2418; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2931 = 4'h3 == io_writeMask ? _GEN_1395 : _GEN_2419; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2932 = 4'h3 == io_writeMask ? _GEN_1396 : _GEN_2420; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2933 = 4'h3 == io_writeMask ? _GEN_1397 : _GEN_2421; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2934 = 4'h3 == io_writeMask ? _GEN_1398 : _GEN_2422; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2935 = 4'h3 == io_writeMask ? _GEN_1399 : _GEN_2423; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2936 = 4'h3 == io_writeMask ? _GEN_1400 : _GEN_2424; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2937 = 4'h3 == io_writeMask ? _GEN_1401 : _GEN_2425; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2938 = 4'h3 == io_writeMask ? _GEN_1402 : _GEN_2426; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2939 = 4'h3 == io_writeMask ? _GEN_1403 : _GEN_2427; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2940 = 4'h3 == io_writeMask ? _GEN_1404 : _GEN_2428; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2941 = 4'h3 == io_writeMask ? _GEN_1405 : _GEN_2429; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2942 = 4'h3 == io_writeMask ? _GEN_1406 : _GEN_2430; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2943 = 4'h3 == io_writeMask ? _GEN_1407 : _GEN_2431; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2944 = 4'h3 == io_writeMask ? _GEN_1408 : _GEN_2432; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2945 = 4'h3 == io_writeMask ? _GEN_1409 : _GEN_2433; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2946 = 4'h3 == io_writeMask ? _GEN_1410 : _GEN_2434; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2947 = 4'h3 == io_writeMask ? _GEN_1411 : _GEN_2435; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2948 = 4'h3 == io_writeMask ? _GEN_1412 : _GEN_2436; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2949 = 4'h3 == io_writeMask ? _GEN_1413 : _GEN_2437; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2950 = 4'h3 == io_writeMask ? _GEN_1414 : _GEN_2438; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2951 = 4'h3 == io_writeMask ? _GEN_1415 : _GEN_2439; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2952 = 4'h3 == io_writeMask ? _GEN_1416 : _GEN_2440; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2953 = 4'h3 == io_writeMask ? _GEN_1417 : _GEN_2441; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2954 = 4'h3 == io_writeMask ? _GEN_1418 : _GEN_2442; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2955 = 4'h3 == io_writeMask ? _GEN_1419 : _GEN_2443; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2956 = 4'h3 == io_writeMask ? _GEN_1420 : _GEN_2444; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2957 = 4'h3 == io_writeMask ? _GEN_1421 : _GEN_2445; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2958 = 4'h3 == io_writeMask ? _GEN_1422 : _GEN_2446; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2959 = 4'h3 == io_writeMask ? _GEN_1423 : _GEN_2447; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2960 = 4'h3 == io_writeMask ? _GEN_1424 : _GEN_2448; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2961 = 4'h3 == io_writeMask ? _GEN_1425 : _GEN_2449; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2962 = 4'h3 == io_writeMask ? _GEN_1426 : _GEN_2450; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2963 = 4'h3 == io_writeMask ? _GEN_1427 : _GEN_2451; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2964 = 4'h3 == io_writeMask ? _GEN_1428 : _GEN_2452; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2965 = 4'h3 == io_writeMask ? _GEN_1429 : _GEN_2453; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2966 = 4'h3 == io_writeMask ? _GEN_1430 : _GEN_2454; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2967 = 4'h3 == io_writeMask ? _GEN_1431 : _GEN_2455; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2968 = 4'h3 == io_writeMask ? _GEN_1432 : _GEN_2456; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2969 = 4'h3 == io_writeMask ? _GEN_1433 : _GEN_2457; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2970 = 4'h3 == io_writeMask ? _GEN_1434 : _GEN_2458; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2971 = 4'h3 == io_writeMask ? _GEN_1435 : _GEN_2459; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2972 = 4'h3 == io_writeMask ? _GEN_1436 : _GEN_2460; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2973 = 4'h3 == io_writeMask ? _GEN_1437 : _GEN_2461; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2974 = 4'h3 == io_writeMask ? _GEN_1438 : _GEN_2462; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2975 = 4'h3 == io_writeMask ? _GEN_1439 : _GEN_2463; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2976 = 4'h3 == io_writeMask ? _GEN_1440 : _GEN_2464; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2977 = 4'h3 == io_writeMask ? _GEN_1441 : _GEN_2465; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2978 = 4'h3 == io_writeMask ? _GEN_1442 : _GEN_2466; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2979 = 4'h3 == io_writeMask ? _GEN_1443 : _GEN_2467; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2980 = 4'h3 == io_writeMask ? _GEN_1444 : _GEN_2468; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2981 = 4'h3 == io_writeMask ? _GEN_1445 : _GEN_2469; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2982 = 4'h3 == io_writeMask ? _GEN_1446 : _GEN_2470; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2983 = 4'h3 == io_writeMask ? _GEN_1447 : _GEN_2471; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2984 = 4'h3 == io_writeMask ? _GEN_1448 : _GEN_2472; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2985 = 4'h3 == io_writeMask ? _GEN_1449 : _GEN_2473; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2986 = 4'h3 == io_writeMask ? _GEN_1450 : _GEN_2474; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2987 = 4'h3 == io_writeMask ? _GEN_1451 : _GEN_2475; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2988 = 4'h3 == io_writeMask ? _GEN_1452 : _GEN_2476; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2989 = 4'h3 == io_writeMask ? _GEN_1453 : _GEN_2477; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2990 = 4'h3 == io_writeMask ? _GEN_1454 : _GEN_2478; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2991 = 4'h3 == io_writeMask ? _GEN_1455 : _GEN_2479; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2992 = 4'h3 == io_writeMask ? _GEN_1456 : _GEN_2480; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2993 = 4'h3 == io_writeMask ? _GEN_1457 : _GEN_2481; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2994 = 4'h3 == io_writeMask ? _GEN_1458 : _GEN_2482; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2995 = 4'h3 == io_writeMask ? _GEN_1459 : _GEN_2483; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2996 = 4'h3 == io_writeMask ? _GEN_1460 : _GEN_2484; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2997 = 4'h3 == io_writeMask ? _GEN_1461 : _GEN_2485; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2998 = 4'h3 == io_writeMask ? _GEN_1462 : _GEN_2486; // @[Cache.scala 133:31]
  wire [31:0] _GEN_2999 = 4'h3 == io_writeMask ? _GEN_1463 : _GEN_2487; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3000 = 4'h3 == io_writeMask ? _GEN_1464 : _GEN_2488; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3001 = 4'h3 == io_writeMask ? _GEN_1465 : _GEN_2489; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3002 = 4'h3 == io_writeMask ? _GEN_1466 : _GEN_2490; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3003 = 4'h3 == io_writeMask ? _GEN_1467 : _GEN_2491; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3004 = 4'h3 == io_writeMask ? _GEN_1468 : _GEN_2492; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3005 = 4'h3 == io_writeMask ? _GEN_1469 : _GEN_2493; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3006 = 4'h3 == io_writeMask ? _GEN_1470 : _GEN_2494; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3007 = 4'h3 == io_writeMask ? _GEN_1471 : _GEN_2495; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3008 = 4'h3 == io_writeMask ? _GEN_1472 : _GEN_2496; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3009 = 4'h3 == io_writeMask ? _GEN_1473 : _GEN_2497; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3010 = 4'h3 == io_writeMask ? _GEN_1474 : _GEN_2498; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3011 = 4'h3 == io_writeMask ? _GEN_1475 : _GEN_2499; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3012 = 4'h3 == io_writeMask ? _GEN_1476 : _GEN_2500; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3013 = 4'h3 == io_writeMask ? _GEN_1477 : _GEN_2501; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3014 = 4'h3 == io_writeMask ? _GEN_1478 : _GEN_2502; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3015 = 4'h3 == io_writeMask ? _GEN_1479 : _GEN_2503; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3016 = 4'h3 == io_writeMask ? _GEN_1480 : _GEN_2504; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3017 = 4'h3 == io_writeMask ? _GEN_1481 : _GEN_2505; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3018 = 4'h3 == io_writeMask ? _GEN_1482 : _GEN_2506; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3019 = 4'h3 == io_writeMask ? _GEN_1483 : _GEN_2507; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3020 = 4'h3 == io_writeMask ? _GEN_1484 : _GEN_2508; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3021 = 4'h3 == io_writeMask ? _GEN_1485 : _GEN_2509; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3022 = 4'h3 == io_writeMask ? _GEN_1486 : _GEN_2510; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3023 = 4'h3 == io_writeMask ? _GEN_1487 : _GEN_2511; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3024 = 4'h3 == io_writeMask ? _GEN_1488 : _GEN_2512; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3025 = 4'h3 == io_writeMask ? _GEN_1489 : _GEN_2513; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3026 = 4'h3 == io_writeMask ? _GEN_1490 : _GEN_2514; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3027 = 4'h3 == io_writeMask ? _GEN_1491 : _GEN_2515; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3028 = 4'h3 == io_writeMask ? _GEN_1492 : _GEN_2516; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3029 = 4'h3 == io_writeMask ? _GEN_1493 : _GEN_2517; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3030 = 4'h3 == io_writeMask ? _GEN_1494 : _GEN_2518; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3031 = 4'h3 == io_writeMask ? _GEN_1495 : _GEN_2519; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3032 = 4'h3 == io_writeMask ? _GEN_1496 : _GEN_2520; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3033 = 4'h3 == io_writeMask ? _GEN_1497 : _GEN_2521; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3034 = 4'h3 == io_writeMask ? _GEN_1498 : _GEN_2522; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3035 = 4'h3 == io_writeMask ? _GEN_1499 : _GEN_2523; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3036 = 4'h3 == io_writeMask ? _GEN_1500 : _GEN_2524; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3037 = 4'h3 == io_writeMask ? _GEN_1501 : _GEN_2525; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3038 = 4'h3 == io_writeMask ? _GEN_1502 : _GEN_2526; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3039 = 4'h3 == io_writeMask ? _GEN_1503 : _GEN_2527; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3040 = 4'h3 == io_writeMask ? _GEN_1504 : _GEN_2528; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3041 = 4'h3 == io_writeMask ? _GEN_1505 : _GEN_2529; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3042 = 4'h3 == io_writeMask ? _GEN_1506 : _GEN_2530; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3043 = 4'h3 == io_writeMask ? _GEN_1507 : _GEN_2531; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3044 = 4'h3 == io_writeMask ? _GEN_1508 : _GEN_2532; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3045 = 4'h3 == io_writeMask ? _GEN_1509 : _GEN_2533; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3046 = 4'h3 == io_writeMask ? _GEN_1510 : _GEN_2534; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3047 = 4'h3 == io_writeMask ? _GEN_1511 : _GEN_2535; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3048 = 4'h3 == io_writeMask ? _GEN_1512 : _GEN_2536; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3049 = 4'h3 == io_writeMask ? _GEN_1513 : _GEN_2537; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3050 = 4'h3 == io_writeMask ? _GEN_1514 : _GEN_2538; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3051 = 4'h3 == io_writeMask ? _GEN_1515 : _GEN_2539; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3052 = 4'h3 == io_writeMask ? _GEN_1516 : _GEN_2540; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3053 = 4'h3 == io_writeMask ? _GEN_1517 : _GEN_2541; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3054 = 4'h3 == io_writeMask ? _GEN_1518 : _GEN_2542; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3055 = 4'h3 == io_writeMask ? _GEN_1519 : _GEN_2543; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3056 = 4'h3 == io_writeMask ? _GEN_1520 : _GEN_2544; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3057 = 4'h3 == io_writeMask ? _GEN_1521 : _GEN_2545; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3058 = 4'h3 == io_writeMask ? _GEN_1522 : _GEN_2546; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3059 = 4'h3 == io_writeMask ? _GEN_1523 : _GEN_2547; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3060 = 4'h3 == io_writeMask ? _GEN_1524 : _GEN_2548; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3061 = 4'h3 == io_writeMask ? _GEN_1525 : _GEN_2549; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3062 = 4'h3 == io_writeMask ? _GEN_1526 : _GEN_2550; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3063 = 4'h3 == io_writeMask ? _GEN_1527 : _GEN_2551; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3064 = 4'h3 == io_writeMask ? _GEN_1528 : _GEN_2552; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3065 = 4'h3 == io_writeMask ? _GEN_1529 : _GEN_2553; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3066 = 4'h3 == io_writeMask ? _GEN_1530 : _GEN_2554; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3067 = 4'h3 == io_writeMask ? _GEN_1531 : _GEN_2555; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3068 = 4'h3 == io_writeMask ? _GEN_1532 : _GEN_2556; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3069 = 4'h3 == io_writeMask ? _GEN_1533 : _GEN_2557; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3070 = 4'h3 == io_writeMask ? _GEN_1534 : _GEN_2558; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3071 = 4'h3 == io_writeMask ? _GEN_1535 : _GEN_2559; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3072 = 4'h3 == io_writeMask ? _GEN_1536 : _GEN_2560; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3073 = 4'h3 == io_writeMask ? _GEN_1537 : _GEN_2561; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3074 = 4'h3 == io_writeMask ? _GEN_1538 : _GEN_2562; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3075 = 4'h3 == io_writeMask ? _GEN_1539 : _GEN_2563; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3076 = 4'h3 == io_writeMask ? _GEN_1540 : _GEN_2564; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3077 = 4'h3 == io_writeMask ? _GEN_1541 : _GEN_2565; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3078 = 4'h3 == io_writeMask ? _GEN_1542 : _GEN_2566; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3079 = 4'h3 == io_writeMask ? _GEN_1543 : _GEN_2567; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3080 = 4'h3 == io_writeMask ? _GEN_1544 : _GEN_2568; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3081 = 4'h3 == io_writeMask ? _GEN_1545 : _GEN_2569; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3082 = 4'h3 == io_writeMask ? _GEN_1546 : _GEN_2570; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3083 = 4'h3 == io_writeMask ? _GEN_1547 : _GEN_2571; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3084 = 4'h3 == io_writeMask ? _GEN_1548 : _GEN_2572; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3085 = 4'h3 == io_writeMask ? _GEN_1549 : _GEN_2573; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3086 = 4'h3 == io_writeMask ? _GEN_1550 : _GEN_2574; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3087 = 4'h3 == io_writeMask ? _GEN_1551 : _GEN_2575; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3088 = 4'h3 == io_writeMask ? _GEN_1552 : _GEN_2576; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3089 = 4'h3 == io_writeMask ? _GEN_1553 : _GEN_2577; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3090 = 4'h3 == io_writeMask ? _GEN_1554 : _GEN_2578; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3091 = 4'h3 == io_writeMask ? _GEN_1555 : _GEN_2579; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3092 = 4'h3 == io_writeMask ? _GEN_1556 : _GEN_2580; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3093 = 4'h3 == io_writeMask ? _GEN_1557 : _GEN_2581; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3094 = 4'h3 == io_writeMask ? _GEN_1558 : _GEN_2582; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3095 = 4'h3 == io_writeMask ? _GEN_1559 : _GEN_2583; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3096 = 4'h3 == io_writeMask ? _GEN_1560 : _GEN_2584; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3097 = 4'h3 == io_writeMask ? _GEN_1561 : _GEN_2585; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3098 = 4'h3 == io_writeMask ? _GEN_1562 : _GEN_2586; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3099 = 4'h3 == io_writeMask ? _GEN_1563 : _GEN_2587; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3100 = 4'h3 == io_writeMask ? _GEN_1564 : _GEN_2588; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3101 = 4'h3 == io_writeMask ? _GEN_1565 : _GEN_2589; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3102 = 4'h3 == io_writeMask ? _GEN_1566 : _GEN_2590; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3103 = 4'h3 == io_writeMask ? _GEN_1567 : _GEN_2591; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3104 = 4'h3 == io_writeMask ? _GEN_1568 : _GEN_2592; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3105 = 4'h3 == io_writeMask ? _GEN_1569 : _GEN_2593; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3106 = 4'h3 == io_writeMask ? _GEN_1570 : _GEN_2594; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3107 = 4'h3 == io_writeMask ? _GEN_1571 : _GEN_2595; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3108 = 4'h3 == io_writeMask ? _GEN_1572 : _GEN_2596; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3109 = 4'h3 == io_writeMask ? _GEN_1573 : _GEN_2597; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3110 = 4'h3 == io_writeMask ? _GEN_1574 : _GEN_2598; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3111 = 4'h3 == io_writeMask ? _GEN_1575 : _GEN_2599; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3112 = 4'h3 == io_writeMask ? _GEN_1576 : _GEN_2600; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3113 = 4'h3 == io_writeMask ? _GEN_1577 : _GEN_2601; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3114 = 4'h3 == io_writeMask ? _GEN_1578 : _GEN_2602; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3115 = 4'h3 == io_writeMask ? _GEN_1579 : _GEN_2603; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3116 = 4'h3 == io_writeMask ? _GEN_1580 : _GEN_2604; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3117 = 4'h3 == io_writeMask ? _GEN_1581 : _GEN_2605; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3118 = 4'h3 == io_writeMask ? _GEN_1582 : _GEN_2606; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3119 = 4'h3 == io_writeMask ? _GEN_1583 : _GEN_2607; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3120 = 4'h3 == io_writeMask ? _GEN_1584 : _GEN_2608; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3121 = 4'h3 == io_writeMask ? _GEN_1585 : _GEN_2609; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3122 = 4'h3 == io_writeMask ? _GEN_1586 : _GEN_2610; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3123 = 4'h3 == io_writeMask ? _GEN_1587 : _GEN_2611; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3124 = 4'h3 == io_writeMask ? _GEN_1588 : _GEN_2612; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3125 = 4'h3 == io_writeMask ? _GEN_1589 : _GEN_2613; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3126 = 4'h3 == io_writeMask ? _GEN_1590 : _GEN_2614; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3127 = 4'h3 == io_writeMask ? _GEN_1591 : _GEN_2615; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3128 = 4'h3 == io_writeMask ? _GEN_1592 : _GEN_2616; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3129 = 4'h3 == io_writeMask ? _GEN_1593 : _GEN_2617; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3130 = 4'h3 == io_writeMask ? _GEN_1594 : _GEN_2618; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3131 = 4'h3 == io_writeMask ? _GEN_1595 : _GEN_2619; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3132 = 4'h3 == io_writeMask ? _GEN_1596 : _GEN_2620; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3133 = 4'h3 == io_writeMask ? _GEN_1597 : _GEN_2621; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3134 = 4'h3 == io_writeMask ? _GEN_1598 : _GEN_2622; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3135 = 4'h3 == io_writeMask ? _GEN_1599 : _GEN_2623; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3136 = 4'h3 == io_writeMask ? _GEN_1600 : _GEN_2624; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3137 = 4'h3 == io_writeMask ? _GEN_1601 : _GEN_2625; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3138 = 4'h3 == io_writeMask ? _GEN_1602 : _GEN_2626; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3139 = 4'h3 == io_writeMask ? _GEN_1603 : _GEN_2627; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3140 = 4'h3 == io_writeMask ? _GEN_1604 : _GEN_2628; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3141 = 4'h3 == io_writeMask ? _GEN_1605 : _GEN_2629; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3142 = 4'h3 == io_writeMask ? _GEN_1606 : _GEN_2630; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3143 = 4'h3 == io_writeMask ? _GEN_1607 : _GEN_2631; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3144 = 4'h3 == io_writeMask ? _GEN_1608 : _GEN_2632; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3145 = 4'h3 == io_writeMask ? _GEN_1609 : _GEN_2633; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3146 = 4'h3 == io_writeMask ? _GEN_1610 : _GEN_2634; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3147 = 4'h3 == io_writeMask ? _GEN_1611 : _GEN_2635; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3148 = 4'h3 == io_writeMask ? _GEN_1612 : _GEN_2636; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3149 = 4'h3 == io_writeMask ? _GEN_1613 : _GEN_2637; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3150 = 4'h3 == io_writeMask ? _GEN_1614 : _GEN_2638; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3151 = 4'h3 == io_writeMask ? _GEN_1615 : _GEN_2639; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3152 = 4'h3 == io_writeMask ? _GEN_1616 : _GEN_2640; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3153 = 4'h3 == io_writeMask ? _GEN_1617 : _GEN_2641; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3154 = 4'h3 == io_writeMask ? _GEN_1618 : _GEN_2642; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3155 = 4'h3 == io_writeMask ? _GEN_1619 : _GEN_2643; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3156 = 4'h3 == io_writeMask ? _GEN_1620 : _GEN_2644; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3157 = 4'h3 == io_writeMask ? _GEN_1621 : _GEN_2645; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3158 = 4'h3 == io_writeMask ? _GEN_1622 : _GEN_2646; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3159 = 4'h3 == io_writeMask ? _GEN_1623 : _GEN_2647; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3160 = 4'h3 == io_writeMask ? _GEN_1624 : _GEN_2648; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3161 = 4'h3 == io_writeMask ? _GEN_1625 : _GEN_2649; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3162 = 4'h3 == io_writeMask ? _GEN_1626 : _GEN_2650; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3163 = 4'h3 == io_writeMask ? _GEN_1627 : _GEN_2651; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3164 = 4'h3 == io_writeMask ? _GEN_1628 : _GEN_2652; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3165 = 4'h3 == io_writeMask ? _GEN_1629 : _GEN_2653; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3166 = 4'h3 == io_writeMask ? _GEN_1630 : _GEN_2654; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3167 = 4'h3 == io_writeMask ? _GEN_1631 : _GEN_2655; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3168 = 4'h3 == io_writeMask ? _GEN_1632 : _GEN_2656; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3169 = 4'h3 == io_writeMask ? _GEN_1633 : _GEN_2657; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3170 = 4'h3 == io_writeMask ? _GEN_1634 : _GEN_2658; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3171 = 4'h3 == io_writeMask ? _GEN_1635 : _GEN_2659; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3172 = 4'h3 == io_writeMask ? _GEN_1636 : _GEN_2660; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3173 = 4'h3 == io_writeMask ? _GEN_1637 : _GEN_2661; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3174 = 4'h3 == io_writeMask ? _GEN_1638 : _GEN_2662; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3175 = 4'h3 == io_writeMask ? _GEN_1639 : _GEN_2663; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3176 = 4'h3 == io_writeMask ? _GEN_1640 : _GEN_2664; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3177 = 4'h3 == io_writeMask ? _GEN_1641 : _GEN_2665; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3178 = 4'h3 == io_writeMask ? _GEN_1642 : _GEN_2666; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3179 = 4'h3 == io_writeMask ? _GEN_1643 : _GEN_2667; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3180 = 4'h3 == io_writeMask ? _GEN_1644 : _GEN_2668; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3181 = 4'h3 == io_writeMask ? _GEN_1645 : _GEN_2669; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3182 = 4'h3 == io_writeMask ? _GEN_1646 : _GEN_2670; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3183 = 4'h3 == io_writeMask ? _GEN_1647 : _GEN_2671; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3184 = 4'h3 == io_writeMask ? _GEN_1648 : _GEN_2672; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3185 = 4'h3 == io_writeMask ? _GEN_1649 : _GEN_2673; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3186 = 4'h3 == io_writeMask ? _GEN_1650 : _GEN_2674; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3187 = 4'h3 == io_writeMask ? _GEN_1651 : _GEN_2675; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3188 = 4'h3 == io_writeMask ? _GEN_1652 : _GEN_2676; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3189 = 4'h3 == io_writeMask ? _GEN_1653 : _GEN_2677; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3190 = 4'h3 == io_writeMask ? _GEN_1654 : _GEN_2678; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3191 = 4'h3 == io_writeMask ? _GEN_1655 : _GEN_2679; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3192 = 4'h3 == io_writeMask ? _GEN_1656 : _GEN_2680; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3193 = 4'h3 == io_writeMask ? _GEN_1657 : _GEN_2681; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3194 = 4'h3 == io_writeMask ? _GEN_1658 : _GEN_2682; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3195 = 4'h3 == io_writeMask ? _GEN_1659 : _GEN_2683; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3196 = 4'h3 == io_writeMask ? _GEN_1660 : _GEN_2684; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3197 = 4'h3 == io_writeMask ? _GEN_1661 : _GEN_2685; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3198 = 4'h3 == io_writeMask ? _GEN_1662 : _GEN_2686; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3199 = 4'h3 == io_writeMask ? _GEN_1663 : _GEN_2687; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3200 = 4'h3 == io_writeMask ? _GEN_1664 : _GEN_2688; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3201 = 4'h3 == io_writeMask ? _GEN_1665 : _GEN_2689; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3202 = 4'h3 == io_writeMask ? _GEN_1666 : _GEN_2690; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3203 = 4'h3 == io_writeMask ? _GEN_1667 : _GEN_2691; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3204 = 4'h3 == io_writeMask ? _GEN_1668 : _GEN_2692; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3205 = 4'h3 == io_writeMask ? _GEN_1669 : _GEN_2693; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3206 = 4'h3 == io_writeMask ? _GEN_1670 : _GEN_2694; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3207 = 4'h3 == io_writeMask ? _GEN_1671 : _GEN_2695; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3208 = 4'h3 == io_writeMask ? _GEN_1672 : _GEN_2696; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3209 = 4'h3 == io_writeMask ? _GEN_1673 : _GEN_2697; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3210 = 4'h3 == io_writeMask ? _GEN_1674 : _GEN_2698; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3211 = 4'h3 == io_writeMask ? _GEN_1675 : _GEN_2699; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3212 = 4'h3 == io_writeMask ? _GEN_1676 : _GEN_2700; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3213 = 4'h3 == io_writeMask ? _GEN_1677 : _GEN_2701; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3214 = 4'h3 == io_writeMask ? _GEN_1678 : _GEN_2702; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3215 = 4'h3 == io_writeMask ? _GEN_1679 : _GEN_2703; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3216 = 4'h3 == io_writeMask ? _GEN_1680 : _GEN_2704; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3217 = 4'h3 == io_writeMask ? _GEN_1681 : _GEN_2705; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3218 = 4'h3 == io_writeMask ? _GEN_1682 : _GEN_2706; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3219 = 4'h3 == io_writeMask ? _GEN_1683 : _GEN_2707; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3220 = 4'h3 == io_writeMask ? _GEN_1684 : _GEN_2708; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3221 = 4'h3 == io_writeMask ? _GEN_1685 : _GEN_2709; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3222 = 4'h3 == io_writeMask ? _GEN_1686 : _GEN_2710; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3223 = 4'h3 == io_writeMask ? _GEN_1687 : _GEN_2711; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3224 = 4'h3 == io_writeMask ? _GEN_1688 : _GEN_2712; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3225 = 4'h3 == io_writeMask ? _GEN_1689 : _GEN_2713; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3226 = 4'h3 == io_writeMask ? _GEN_1690 : _GEN_2714; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3227 = 4'h3 == io_writeMask ? _GEN_1691 : _GEN_2715; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3228 = 4'h3 == io_writeMask ? _GEN_1692 : _GEN_2716; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3229 = 4'h3 == io_writeMask ? _GEN_1693 : _GEN_2717; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3230 = 4'h3 == io_writeMask ? _GEN_1694 : _GEN_2718; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3231 = 4'h3 == io_writeMask ? _GEN_1695 : _GEN_2719; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3232 = 4'h3 == io_writeMask ? _GEN_1696 : _GEN_2720; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3233 = 4'h3 == io_writeMask ? _GEN_1697 : _GEN_2721; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3234 = 4'h3 == io_writeMask ? _GEN_1698 : _GEN_2722; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3235 = 4'h3 == io_writeMask ? _GEN_1699 : _GEN_2723; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3236 = 4'h3 == io_writeMask ? _GEN_1700 : _GEN_2724; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3237 = 4'h3 == io_writeMask ? _GEN_1701 : _GEN_2725; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3238 = 4'h3 == io_writeMask ? _GEN_1702 : _GEN_2726; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3239 = 4'h3 == io_writeMask ? _GEN_1703 : _GEN_2727; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3240 = 4'h3 == io_writeMask ? _GEN_1704 : _GEN_2728; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3241 = 4'h3 == io_writeMask ? _GEN_1705 : _GEN_2729; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3242 = 4'h3 == io_writeMask ? _GEN_1706 : _GEN_2730; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3243 = 4'h3 == io_writeMask ? _GEN_1707 : _GEN_2731; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3244 = 4'h3 == io_writeMask ? _GEN_1708 : _GEN_2732; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3245 = 4'h3 == io_writeMask ? _GEN_1709 : _GEN_2733; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3246 = 4'h3 == io_writeMask ? _GEN_1710 : _GEN_2734; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3247 = 4'h3 == io_writeMask ? _GEN_1711 : _GEN_2735; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3248 = 4'h3 == io_writeMask ? _GEN_1712 : _GEN_2736; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3249 = 4'h3 == io_writeMask ? _GEN_1713 : _GEN_2737; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3250 = 4'h3 == io_writeMask ? _GEN_1714 : _GEN_2738; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3251 = 4'h1 == io_writeMask ? _GEN_691 : _GEN_2739; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3252 = 4'h1 == io_writeMask ? _GEN_692 : _GEN_2740; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3253 = 4'h1 == io_writeMask ? _GEN_693 : _GEN_2741; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3254 = 4'h1 == io_writeMask ? _GEN_694 : _GEN_2742; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3255 = 4'h1 == io_writeMask ? _GEN_695 : _GEN_2743; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3256 = 4'h1 == io_writeMask ? _GEN_696 : _GEN_2744; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3257 = 4'h1 == io_writeMask ? _GEN_697 : _GEN_2745; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3258 = 4'h1 == io_writeMask ? _GEN_698 : _GEN_2746; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3259 = 4'h1 == io_writeMask ? _GEN_699 : _GEN_2747; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3260 = 4'h1 == io_writeMask ? _GEN_700 : _GEN_2748; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3261 = 4'h1 == io_writeMask ? _GEN_701 : _GEN_2749; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3262 = 4'h1 == io_writeMask ? _GEN_702 : _GEN_2750; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3263 = 4'h1 == io_writeMask ? _GEN_703 : _GEN_2751; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3264 = 4'h1 == io_writeMask ? _GEN_704 : _GEN_2752; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3265 = 4'h1 == io_writeMask ? _GEN_705 : _GEN_2753; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3266 = 4'h1 == io_writeMask ? _GEN_706 : _GEN_2754; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3267 = 4'h1 == io_writeMask ? _GEN_707 : _GEN_2755; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3268 = 4'h1 == io_writeMask ? _GEN_708 : _GEN_2756; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3269 = 4'h1 == io_writeMask ? _GEN_709 : _GEN_2757; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3270 = 4'h1 == io_writeMask ? _GEN_710 : _GEN_2758; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3271 = 4'h1 == io_writeMask ? _GEN_711 : _GEN_2759; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3272 = 4'h1 == io_writeMask ? _GEN_712 : _GEN_2760; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3273 = 4'h1 == io_writeMask ? _GEN_713 : _GEN_2761; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3274 = 4'h1 == io_writeMask ? _GEN_714 : _GEN_2762; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3275 = 4'h1 == io_writeMask ? _GEN_715 : _GEN_2763; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3276 = 4'h1 == io_writeMask ? _GEN_716 : _GEN_2764; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3277 = 4'h1 == io_writeMask ? _GEN_717 : _GEN_2765; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3278 = 4'h1 == io_writeMask ? _GEN_718 : _GEN_2766; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3279 = 4'h1 == io_writeMask ? _GEN_719 : _GEN_2767; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3280 = 4'h1 == io_writeMask ? _GEN_720 : _GEN_2768; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3281 = 4'h1 == io_writeMask ? _GEN_721 : _GEN_2769; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3282 = 4'h1 == io_writeMask ? _GEN_722 : _GEN_2770; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3283 = 4'h1 == io_writeMask ? _GEN_723 : _GEN_2771; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3284 = 4'h1 == io_writeMask ? _GEN_724 : _GEN_2772; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3285 = 4'h1 == io_writeMask ? _GEN_725 : _GEN_2773; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3286 = 4'h1 == io_writeMask ? _GEN_726 : _GEN_2774; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3287 = 4'h1 == io_writeMask ? _GEN_727 : _GEN_2775; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3288 = 4'h1 == io_writeMask ? _GEN_728 : _GEN_2776; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3289 = 4'h1 == io_writeMask ? _GEN_729 : _GEN_2777; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3290 = 4'h1 == io_writeMask ? _GEN_730 : _GEN_2778; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3291 = 4'h1 == io_writeMask ? _GEN_731 : _GEN_2779; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3292 = 4'h1 == io_writeMask ? _GEN_732 : _GEN_2780; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3293 = 4'h1 == io_writeMask ? _GEN_733 : _GEN_2781; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3294 = 4'h1 == io_writeMask ? _GEN_734 : _GEN_2782; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3295 = 4'h1 == io_writeMask ? _GEN_735 : _GEN_2783; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3296 = 4'h1 == io_writeMask ? _GEN_736 : _GEN_2784; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3297 = 4'h1 == io_writeMask ? _GEN_737 : _GEN_2785; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3298 = 4'h1 == io_writeMask ? _GEN_738 : _GEN_2786; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3299 = 4'h1 == io_writeMask ? _GEN_739 : _GEN_2787; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3300 = 4'h1 == io_writeMask ? _GEN_740 : _GEN_2788; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3301 = 4'h1 == io_writeMask ? _GEN_741 : _GEN_2789; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3302 = 4'h1 == io_writeMask ? _GEN_742 : _GEN_2790; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3303 = 4'h1 == io_writeMask ? _GEN_743 : _GEN_2791; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3304 = 4'h1 == io_writeMask ? _GEN_744 : _GEN_2792; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3305 = 4'h1 == io_writeMask ? _GEN_745 : _GEN_2793; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3306 = 4'h1 == io_writeMask ? _GEN_746 : _GEN_2794; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3307 = 4'h1 == io_writeMask ? _GEN_747 : _GEN_2795; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3308 = 4'h1 == io_writeMask ? _GEN_748 : _GEN_2796; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3309 = 4'h1 == io_writeMask ? _GEN_749 : _GEN_2797; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3310 = 4'h1 == io_writeMask ? _GEN_750 : _GEN_2798; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3311 = 4'h1 == io_writeMask ? _GEN_751 : _GEN_2799; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3312 = 4'h1 == io_writeMask ? _GEN_752 : _GEN_2800; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3313 = 4'h1 == io_writeMask ? _GEN_753 : _GEN_2801; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3314 = 4'h1 == io_writeMask ? _GEN_754 : _GEN_2802; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3315 = 4'h1 == io_writeMask ? _GEN_755 : _GEN_2803; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3316 = 4'h1 == io_writeMask ? _GEN_756 : _GEN_2804; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3317 = 4'h1 == io_writeMask ? _GEN_757 : _GEN_2805; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3318 = 4'h1 == io_writeMask ? _GEN_758 : _GEN_2806; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3319 = 4'h1 == io_writeMask ? _GEN_759 : _GEN_2807; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3320 = 4'h1 == io_writeMask ? _GEN_760 : _GEN_2808; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3321 = 4'h1 == io_writeMask ? _GEN_761 : _GEN_2809; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3322 = 4'h1 == io_writeMask ? _GEN_762 : _GEN_2810; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3323 = 4'h1 == io_writeMask ? _GEN_763 : _GEN_2811; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3324 = 4'h1 == io_writeMask ? _GEN_764 : _GEN_2812; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3325 = 4'h1 == io_writeMask ? _GEN_765 : _GEN_2813; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3326 = 4'h1 == io_writeMask ? _GEN_766 : _GEN_2814; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3327 = 4'h1 == io_writeMask ? _GEN_767 : _GEN_2815; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3328 = 4'h1 == io_writeMask ? _GEN_768 : _GEN_2816; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3329 = 4'h1 == io_writeMask ? _GEN_769 : _GEN_2817; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3330 = 4'h1 == io_writeMask ? _GEN_770 : _GEN_2818; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3331 = 4'h1 == io_writeMask ? _GEN_771 : _GEN_2819; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3332 = 4'h1 == io_writeMask ? _GEN_772 : _GEN_2820; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3333 = 4'h1 == io_writeMask ? _GEN_773 : _GEN_2821; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3334 = 4'h1 == io_writeMask ? _GEN_774 : _GEN_2822; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3335 = 4'h1 == io_writeMask ? _GEN_775 : _GEN_2823; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3336 = 4'h1 == io_writeMask ? _GEN_776 : _GEN_2824; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3337 = 4'h1 == io_writeMask ? _GEN_777 : _GEN_2825; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3338 = 4'h1 == io_writeMask ? _GEN_778 : _GEN_2826; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3339 = 4'h1 == io_writeMask ? _GEN_779 : _GEN_2827; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3340 = 4'h1 == io_writeMask ? _GEN_780 : _GEN_2828; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3341 = 4'h1 == io_writeMask ? _GEN_781 : _GEN_2829; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3342 = 4'h1 == io_writeMask ? _GEN_782 : _GEN_2830; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3343 = 4'h1 == io_writeMask ? _GEN_783 : _GEN_2831; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3344 = 4'h1 == io_writeMask ? _GEN_784 : _GEN_2832; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3345 = 4'h1 == io_writeMask ? _GEN_785 : _GEN_2833; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3346 = 4'h1 == io_writeMask ? _GEN_786 : _GEN_2834; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3347 = 4'h1 == io_writeMask ? _GEN_787 : _GEN_2835; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3348 = 4'h1 == io_writeMask ? _GEN_788 : _GEN_2836; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3349 = 4'h1 == io_writeMask ? _GEN_789 : _GEN_2837; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3350 = 4'h1 == io_writeMask ? _GEN_790 : _GEN_2838; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3351 = 4'h1 == io_writeMask ? _GEN_791 : _GEN_2839; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3352 = 4'h1 == io_writeMask ? _GEN_792 : _GEN_2840; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3353 = 4'h1 == io_writeMask ? _GEN_793 : _GEN_2841; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3354 = 4'h1 == io_writeMask ? _GEN_794 : _GEN_2842; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3355 = 4'h1 == io_writeMask ? _GEN_795 : _GEN_2843; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3356 = 4'h1 == io_writeMask ? _GEN_796 : _GEN_2844; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3357 = 4'h1 == io_writeMask ? _GEN_797 : _GEN_2845; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3358 = 4'h1 == io_writeMask ? _GEN_798 : _GEN_2846; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3359 = 4'h1 == io_writeMask ? _GEN_799 : _GEN_2847; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3360 = 4'h1 == io_writeMask ? _GEN_800 : _GEN_2848; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3361 = 4'h1 == io_writeMask ? _GEN_801 : _GEN_2849; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3362 = 4'h1 == io_writeMask ? _GEN_802 : _GEN_2850; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3363 = 4'h1 == io_writeMask ? _GEN_803 : _GEN_2851; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3364 = 4'h1 == io_writeMask ? _GEN_804 : _GEN_2852; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3365 = 4'h1 == io_writeMask ? _GEN_805 : _GEN_2853; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3366 = 4'h1 == io_writeMask ? _GEN_806 : _GEN_2854; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3367 = 4'h1 == io_writeMask ? _GEN_807 : _GEN_2855; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3368 = 4'h1 == io_writeMask ? _GEN_808 : _GEN_2856; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3369 = 4'h1 == io_writeMask ? _GEN_809 : _GEN_2857; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3370 = 4'h1 == io_writeMask ? _GEN_810 : _GEN_2858; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3371 = 4'h1 == io_writeMask ? _GEN_811 : _GEN_2859; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3372 = 4'h1 == io_writeMask ? _GEN_812 : _GEN_2860; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3373 = 4'h1 == io_writeMask ? _GEN_813 : _GEN_2861; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3374 = 4'h1 == io_writeMask ? _GEN_814 : _GEN_2862; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3375 = 4'h1 == io_writeMask ? _GEN_815 : _GEN_2863; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3376 = 4'h1 == io_writeMask ? _GEN_816 : _GEN_2864; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3377 = 4'h1 == io_writeMask ? _GEN_817 : _GEN_2865; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3378 = 4'h1 == io_writeMask ? _GEN_818 : _GEN_2866; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3379 = 4'h1 == io_writeMask ? _GEN_819 : _GEN_2867; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3380 = 4'h1 == io_writeMask ? _GEN_820 : _GEN_2868; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3381 = 4'h1 == io_writeMask ? _GEN_821 : _GEN_2869; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3382 = 4'h1 == io_writeMask ? _GEN_822 : _GEN_2870; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3383 = 4'h1 == io_writeMask ? _GEN_823 : _GEN_2871; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3384 = 4'h1 == io_writeMask ? _GEN_824 : _GEN_2872; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3385 = 4'h1 == io_writeMask ? _GEN_825 : _GEN_2873; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3386 = 4'h1 == io_writeMask ? _GEN_826 : _GEN_2874; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3387 = 4'h1 == io_writeMask ? _GEN_827 : _GEN_2875; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3388 = 4'h1 == io_writeMask ? _GEN_828 : _GEN_2876; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3389 = 4'h1 == io_writeMask ? _GEN_829 : _GEN_2877; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3390 = 4'h1 == io_writeMask ? _GEN_830 : _GEN_2878; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3391 = 4'h1 == io_writeMask ? _GEN_831 : _GEN_2879; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3392 = 4'h1 == io_writeMask ? _GEN_832 : _GEN_2880; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3393 = 4'h1 == io_writeMask ? _GEN_833 : _GEN_2881; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3394 = 4'h1 == io_writeMask ? _GEN_834 : _GEN_2882; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3395 = 4'h1 == io_writeMask ? _GEN_835 : _GEN_2883; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3396 = 4'h1 == io_writeMask ? _GEN_836 : _GEN_2884; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3397 = 4'h1 == io_writeMask ? _GEN_837 : _GEN_2885; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3398 = 4'h1 == io_writeMask ? _GEN_838 : _GEN_2886; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3399 = 4'h1 == io_writeMask ? _GEN_839 : _GEN_2887; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3400 = 4'h1 == io_writeMask ? _GEN_840 : _GEN_2888; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3401 = 4'h1 == io_writeMask ? _GEN_841 : _GEN_2889; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3402 = 4'h1 == io_writeMask ? _GEN_842 : _GEN_2890; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3403 = 4'h1 == io_writeMask ? _GEN_843 : _GEN_2891; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3404 = 4'h1 == io_writeMask ? _GEN_844 : _GEN_2892; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3405 = 4'h1 == io_writeMask ? _GEN_845 : _GEN_2893; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3406 = 4'h1 == io_writeMask ? _GEN_846 : _GEN_2894; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3407 = 4'h1 == io_writeMask ? _GEN_847 : _GEN_2895; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3408 = 4'h1 == io_writeMask ? _GEN_848 : _GEN_2896; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3409 = 4'h1 == io_writeMask ? _GEN_849 : _GEN_2897; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3410 = 4'h1 == io_writeMask ? _GEN_850 : _GEN_2898; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3411 = 4'h1 == io_writeMask ? _GEN_851 : _GEN_2899; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3412 = 4'h1 == io_writeMask ? _GEN_852 : _GEN_2900; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3413 = 4'h1 == io_writeMask ? _GEN_853 : _GEN_2901; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3414 = 4'h1 == io_writeMask ? _GEN_854 : _GEN_2902; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3415 = 4'h1 == io_writeMask ? _GEN_855 : _GEN_2903; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3416 = 4'h1 == io_writeMask ? _GEN_856 : _GEN_2904; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3417 = 4'h1 == io_writeMask ? _GEN_857 : _GEN_2905; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3418 = 4'h1 == io_writeMask ? _GEN_858 : _GEN_2906; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3419 = 4'h1 == io_writeMask ? _GEN_859 : _GEN_2907; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3420 = 4'h1 == io_writeMask ? _GEN_860 : _GEN_2908; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3421 = 4'h1 == io_writeMask ? _GEN_861 : _GEN_2909; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3422 = 4'h1 == io_writeMask ? _GEN_862 : _GEN_2910; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3423 = 4'h1 == io_writeMask ? _GEN_863 : _GEN_2911; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3424 = 4'h1 == io_writeMask ? _GEN_864 : _GEN_2912; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3425 = 4'h1 == io_writeMask ? _GEN_865 : _GEN_2913; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3426 = 4'h1 == io_writeMask ? _GEN_866 : _GEN_2914; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3427 = 4'h1 == io_writeMask ? _GEN_867 : _GEN_2915; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3428 = 4'h1 == io_writeMask ? _GEN_868 : _GEN_2916; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3429 = 4'h1 == io_writeMask ? _GEN_869 : _GEN_2917; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3430 = 4'h1 == io_writeMask ? _GEN_870 : _GEN_2918; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3431 = 4'h1 == io_writeMask ? _GEN_871 : _GEN_2919; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3432 = 4'h1 == io_writeMask ? _GEN_872 : _GEN_2920; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3433 = 4'h1 == io_writeMask ? _GEN_873 : _GEN_2921; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3434 = 4'h1 == io_writeMask ? _GEN_874 : _GEN_2922; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3435 = 4'h1 == io_writeMask ? _GEN_875 : _GEN_2923; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3436 = 4'h1 == io_writeMask ? _GEN_876 : _GEN_2924; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3437 = 4'h1 == io_writeMask ? _GEN_877 : _GEN_2925; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3438 = 4'h1 == io_writeMask ? _GEN_878 : _GEN_2926; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3439 = 4'h1 == io_writeMask ? _GEN_879 : _GEN_2927; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3440 = 4'h1 == io_writeMask ? _GEN_880 : _GEN_2928; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3441 = 4'h1 == io_writeMask ? _GEN_881 : _GEN_2929; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3442 = 4'h1 == io_writeMask ? _GEN_882 : _GEN_2930; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3443 = 4'h1 == io_writeMask ? _GEN_883 : _GEN_2931; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3444 = 4'h1 == io_writeMask ? _GEN_884 : _GEN_2932; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3445 = 4'h1 == io_writeMask ? _GEN_885 : _GEN_2933; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3446 = 4'h1 == io_writeMask ? _GEN_886 : _GEN_2934; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3447 = 4'h1 == io_writeMask ? _GEN_887 : _GEN_2935; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3448 = 4'h1 == io_writeMask ? _GEN_888 : _GEN_2936; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3449 = 4'h1 == io_writeMask ? _GEN_889 : _GEN_2937; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3450 = 4'h1 == io_writeMask ? _GEN_890 : _GEN_2938; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3451 = 4'h1 == io_writeMask ? _GEN_891 : _GEN_2939; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3452 = 4'h1 == io_writeMask ? _GEN_892 : _GEN_2940; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3453 = 4'h1 == io_writeMask ? _GEN_893 : _GEN_2941; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3454 = 4'h1 == io_writeMask ? _GEN_894 : _GEN_2942; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3455 = 4'h1 == io_writeMask ? _GEN_895 : _GEN_2943; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3456 = 4'h1 == io_writeMask ? _GEN_896 : _GEN_2944; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3457 = 4'h1 == io_writeMask ? _GEN_897 : _GEN_2945; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3458 = 4'h1 == io_writeMask ? _GEN_898 : _GEN_2946; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3459 = 4'h1 == io_writeMask ? _GEN_899 : _GEN_2947; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3460 = 4'h1 == io_writeMask ? _GEN_900 : _GEN_2948; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3461 = 4'h1 == io_writeMask ? _GEN_901 : _GEN_2949; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3462 = 4'h1 == io_writeMask ? _GEN_902 : _GEN_2950; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3463 = 4'h1 == io_writeMask ? _GEN_903 : _GEN_2951; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3464 = 4'h1 == io_writeMask ? _GEN_904 : _GEN_2952; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3465 = 4'h1 == io_writeMask ? _GEN_905 : _GEN_2953; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3466 = 4'h1 == io_writeMask ? _GEN_906 : _GEN_2954; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3467 = 4'h1 == io_writeMask ? _GEN_907 : _GEN_2955; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3468 = 4'h1 == io_writeMask ? _GEN_908 : _GEN_2956; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3469 = 4'h1 == io_writeMask ? _GEN_909 : _GEN_2957; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3470 = 4'h1 == io_writeMask ? _GEN_910 : _GEN_2958; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3471 = 4'h1 == io_writeMask ? _GEN_911 : _GEN_2959; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3472 = 4'h1 == io_writeMask ? _GEN_912 : _GEN_2960; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3473 = 4'h1 == io_writeMask ? _GEN_913 : _GEN_2961; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3474 = 4'h1 == io_writeMask ? _GEN_914 : _GEN_2962; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3475 = 4'h1 == io_writeMask ? _GEN_915 : _GEN_2963; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3476 = 4'h1 == io_writeMask ? _GEN_916 : _GEN_2964; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3477 = 4'h1 == io_writeMask ? _GEN_917 : _GEN_2965; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3478 = 4'h1 == io_writeMask ? _GEN_918 : _GEN_2966; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3479 = 4'h1 == io_writeMask ? _GEN_919 : _GEN_2967; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3480 = 4'h1 == io_writeMask ? _GEN_920 : _GEN_2968; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3481 = 4'h1 == io_writeMask ? _GEN_921 : _GEN_2969; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3482 = 4'h1 == io_writeMask ? _GEN_922 : _GEN_2970; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3483 = 4'h1 == io_writeMask ? _GEN_923 : _GEN_2971; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3484 = 4'h1 == io_writeMask ? _GEN_924 : _GEN_2972; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3485 = 4'h1 == io_writeMask ? _GEN_925 : _GEN_2973; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3486 = 4'h1 == io_writeMask ? _GEN_926 : _GEN_2974; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3487 = 4'h1 == io_writeMask ? _GEN_927 : _GEN_2975; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3488 = 4'h1 == io_writeMask ? _GEN_928 : _GEN_2976; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3489 = 4'h1 == io_writeMask ? _GEN_929 : _GEN_2977; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3490 = 4'h1 == io_writeMask ? _GEN_930 : _GEN_2978; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3491 = 4'h1 == io_writeMask ? _GEN_931 : _GEN_2979; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3492 = 4'h1 == io_writeMask ? _GEN_932 : _GEN_2980; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3493 = 4'h1 == io_writeMask ? _GEN_933 : _GEN_2981; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3494 = 4'h1 == io_writeMask ? _GEN_934 : _GEN_2982; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3495 = 4'h1 == io_writeMask ? _GEN_935 : _GEN_2983; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3496 = 4'h1 == io_writeMask ? _GEN_936 : _GEN_2984; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3497 = 4'h1 == io_writeMask ? _GEN_937 : _GEN_2985; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3498 = 4'h1 == io_writeMask ? _GEN_938 : _GEN_2986; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3499 = 4'h1 == io_writeMask ? _GEN_939 : _GEN_2987; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3500 = 4'h1 == io_writeMask ? _GEN_940 : _GEN_2988; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3501 = 4'h1 == io_writeMask ? _GEN_941 : _GEN_2989; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3502 = 4'h1 == io_writeMask ? _GEN_942 : _GEN_2990; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3503 = 4'h1 == io_writeMask ? _GEN_943 : _GEN_2991; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3504 = 4'h1 == io_writeMask ? _GEN_944 : _GEN_2992; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3505 = 4'h1 == io_writeMask ? _GEN_945 : _GEN_2993; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3506 = 4'h1 == io_writeMask ? _GEN_946 : _GEN_2994; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3507 = 4'h1 == io_writeMask ? _GEN_947 : _GEN_2995; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3508 = 4'h1 == io_writeMask ? _GEN_948 : _GEN_2996; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3509 = 4'h1 == io_writeMask ? _GEN_949 : _GEN_2997; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3510 = 4'h1 == io_writeMask ? _GEN_950 : _GEN_2998; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3511 = 4'h1 == io_writeMask ? _GEN_951 : _GEN_2999; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3512 = 4'h1 == io_writeMask ? _GEN_952 : _GEN_3000; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3513 = 4'h1 == io_writeMask ? _GEN_953 : _GEN_3001; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3514 = 4'h1 == io_writeMask ? _GEN_954 : _GEN_3002; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3515 = 4'h1 == io_writeMask ? _GEN_955 : _GEN_3003; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3516 = 4'h1 == io_writeMask ? _GEN_956 : _GEN_3004; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3517 = 4'h1 == io_writeMask ? _GEN_957 : _GEN_3005; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3518 = 4'h1 == io_writeMask ? _GEN_958 : _GEN_3006; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3519 = 4'h1 == io_writeMask ? _GEN_959 : _GEN_3007; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3520 = 4'h1 == io_writeMask ? _GEN_960 : _GEN_3008; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3521 = 4'h1 == io_writeMask ? _GEN_961 : _GEN_3009; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3522 = 4'h1 == io_writeMask ? _GEN_962 : _GEN_3010; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3523 = 4'h1 == io_writeMask ? _GEN_963 : _GEN_3011; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3524 = 4'h1 == io_writeMask ? _GEN_964 : _GEN_3012; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3525 = 4'h1 == io_writeMask ? _GEN_965 : _GEN_3013; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3526 = 4'h1 == io_writeMask ? _GEN_966 : _GEN_3014; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3527 = 4'h1 == io_writeMask ? _GEN_967 : _GEN_3015; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3528 = 4'h1 == io_writeMask ? _GEN_968 : _GEN_3016; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3529 = 4'h1 == io_writeMask ? _GEN_969 : _GEN_3017; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3530 = 4'h1 == io_writeMask ? _GEN_970 : _GEN_3018; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3531 = 4'h1 == io_writeMask ? _GEN_971 : _GEN_3019; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3532 = 4'h1 == io_writeMask ? _GEN_972 : _GEN_3020; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3533 = 4'h1 == io_writeMask ? _GEN_973 : _GEN_3021; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3534 = 4'h1 == io_writeMask ? _GEN_974 : _GEN_3022; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3535 = 4'h1 == io_writeMask ? _GEN_975 : _GEN_3023; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3536 = 4'h1 == io_writeMask ? _GEN_976 : _GEN_3024; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3537 = 4'h1 == io_writeMask ? _GEN_977 : _GEN_3025; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3538 = 4'h1 == io_writeMask ? _GEN_978 : _GEN_3026; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3539 = 4'h1 == io_writeMask ? _GEN_979 : _GEN_3027; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3540 = 4'h1 == io_writeMask ? _GEN_980 : _GEN_3028; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3541 = 4'h1 == io_writeMask ? _GEN_981 : _GEN_3029; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3542 = 4'h1 == io_writeMask ? _GEN_982 : _GEN_3030; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3543 = 4'h1 == io_writeMask ? _GEN_983 : _GEN_3031; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3544 = 4'h1 == io_writeMask ? _GEN_984 : _GEN_3032; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3545 = 4'h1 == io_writeMask ? _GEN_985 : _GEN_3033; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3546 = 4'h1 == io_writeMask ? _GEN_986 : _GEN_3034; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3547 = 4'h1 == io_writeMask ? _GEN_987 : _GEN_3035; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3548 = 4'h1 == io_writeMask ? _GEN_988 : _GEN_3036; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3549 = 4'h1 == io_writeMask ? _GEN_989 : _GEN_3037; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3550 = 4'h1 == io_writeMask ? _GEN_990 : _GEN_3038; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3551 = 4'h1 == io_writeMask ? _GEN_991 : _GEN_3039; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3552 = 4'h1 == io_writeMask ? _GEN_992 : _GEN_3040; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3553 = 4'h1 == io_writeMask ? _GEN_993 : _GEN_3041; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3554 = 4'h1 == io_writeMask ? _GEN_994 : _GEN_3042; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3555 = 4'h1 == io_writeMask ? _GEN_995 : _GEN_3043; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3556 = 4'h1 == io_writeMask ? _GEN_996 : _GEN_3044; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3557 = 4'h1 == io_writeMask ? _GEN_997 : _GEN_3045; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3558 = 4'h1 == io_writeMask ? _GEN_998 : _GEN_3046; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3559 = 4'h1 == io_writeMask ? _GEN_999 : _GEN_3047; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3560 = 4'h1 == io_writeMask ? _GEN_1000 : _GEN_3048; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3561 = 4'h1 == io_writeMask ? _GEN_1001 : _GEN_3049; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3562 = 4'h1 == io_writeMask ? _GEN_1002 : _GEN_3050; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3563 = 4'h1 == io_writeMask ? _GEN_1003 : _GEN_3051; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3564 = 4'h1 == io_writeMask ? _GEN_1004 : _GEN_3052; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3565 = 4'h1 == io_writeMask ? _GEN_1005 : _GEN_3053; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3566 = 4'h1 == io_writeMask ? _GEN_1006 : _GEN_3054; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3567 = 4'h1 == io_writeMask ? _GEN_1007 : _GEN_3055; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3568 = 4'h1 == io_writeMask ? _GEN_1008 : _GEN_3056; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3569 = 4'h1 == io_writeMask ? _GEN_1009 : _GEN_3057; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3570 = 4'h1 == io_writeMask ? _GEN_1010 : _GEN_3058; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3571 = 4'h1 == io_writeMask ? _GEN_1011 : _GEN_3059; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3572 = 4'h1 == io_writeMask ? _GEN_1012 : _GEN_3060; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3573 = 4'h1 == io_writeMask ? _GEN_1013 : _GEN_3061; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3574 = 4'h1 == io_writeMask ? _GEN_1014 : _GEN_3062; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3575 = 4'h1 == io_writeMask ? _GEN_1015 : _GEN_3063; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3576 = 4'h1 == io_writeMask ? _GEN_1016 : _GEN_3064; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3577 = 4'h1 == io_writeMask ? _GEN_1017 : _GEN_3065; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3578 = 4'h1 == io_writeMask ? _GEN_1018 : _GEN_3066; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3579 = 4'h1 == io_writeMask ? _GEN_1019 : _GEN_3067; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3580 = 4'h1 == io_writeMask ? _GEN_1020 : _GEN_3068; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3581 = 4'h1 == io_writeMask ? _GEN_1021 : _GEN_3069; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3582 = 4'h1 == io_writeMask ? _GEN_1022 : _GEN_3070; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3583 = 4'h1 == io_writeMask ? _GEN_1023 : _GEN_3071; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3584 = 4'h1 == io_writeMask ? _GEN_1024 : _GEN_3072; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3585 = 4'h1 == io_writeMask ? _GEN_1025 : _GEN_3073; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3586 = 4'h1 == io_writeMask ? _GEN_1026 : _GEN_3074; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3587 = 4'h1 == io_writeMask ? _GEN_1027 : _GEN_3075; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3588 = 4'h1 == io_writeMask ? _GEN_1028 : _GEN_3076; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3589 = 4'h1 == io_writeMask ? _GEN_1029 : _GEN_3077; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3590 = 4'h1 == io_writeMask ? _GEN_1030 : _GEN_3078; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3591 = 4'h1 == io_writeMask ? _GEN_1031 : _GEN_3079; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3592 = 4'h1 == io_writeMask ? _GEN_1032 : _GEN_3080; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3593 = 4'h1 == io_writeMask ? _GEN_1033 : _GEN_3081; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3594 = 4'h1 == io_writeMask ? _GEN_1034 : _GEN_3082; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3595 = 4'h1 == io_writeMask ? _GEN_1035 : _GEN_3083; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3596 = 4'h1 == io_writeMask ? _GEN_1036 : _GEN_3084; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3597 = 4'h1 == io_writeMask ? _GEN_1037 : _GEN_3085; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3598 = 4'h1 == io_writeMask ? _GEN_1038 : _GEN_3086; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3599 = 4'h1 == io_writeMask ? _GEN_1039 : _GEN_3087; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3600 = 4'h1 == io_writeMask ? _GEN_1040 : _GEN_3088; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3601 = 4'h1 == io_writeMask ? _GEN_1041 : _GEN_3089; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3602 = 4'h1 == io_writeMask ? _GEN_1042 : _GEN_3090; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3603 = 4'h1 == io_writeMask ? _GEN_1043 : _GEN_3091; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3604 = 4'h1 == io_writeMask ? _GEN_1044 : _GEN_3092; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3605 = 4'h1 == io_writeMask ? _GEN_1045 : _GEN_3093; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3606 = 4'h1 == io_writeMask ? _GEN_1046 : _GEN_3094; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3607 = 4'h1 == io_writeMask ? _GEN_1047 : _GEN_3095; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3608 = 4'h1 == io_writeMask ? _GEN_1048 : _GEN_3096; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3609 = 4'h1 == io_writeMask ? _GEN_1049 : _GEN_3097; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3610 = 4'h1 == io_writeMask ? _GEN_1050 : _GEN_3098; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3611 = 4'h1 == io_writeMask ? _GEN_1051 : _GEN_3099; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3612 = 4'h1 == io_writeMask ? _GEN_1052 : _GEN_3100; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3613 = 4'h1 == io_writeMask ? _GEN_1053 : _GEN_3101; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3614 = 4'h1 == io_writeMask ? _GEN_1054 : _GEN_3102; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3615 = 4'h1 == io_writeMask ? _GEN_1055 : _GEN_3103; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3616 = 4'h1 == io_writeMask ? _GEN_1056 : _GEN_3104; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3617 = 4'h1 == io_writeMask ? _GEN_1057 : _GEN_3105; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3618 = 4'h1 == io_writeMask ? _GEN_1058 : _GEN_3106; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3619 = 4'h1 == io_writeMask ? _GEN_1059 : _GEN_3107; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3620 = 4'h1 == io_writeMask ? _GEN_1060 : _GEN_3108; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3621 = 4'h1 == io_writeMask ? _GEN_1061 : _GEN_3109; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3622 = 4'h1 == io_writeMask ? _GEN_1062 : _GEN_3110; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3623 = 4'h1 == io_writeMask ? _GEN_1063 : _GEN_3111; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3624 = 4'h1 == io_writeMask ? _GEN_1064 : _GEN_3112; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3625 = 4'h1 == io_writeMask ? _GEN_1065 : _GEN_3113; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3626 = 4'h1 == io_writeMask ? _GEN_1066 : _GEN_3114; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3627 = 4'h1 == io_writeMask ? _GEN_1067 : _GEN_3115; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3628 = 4'h1 == io_writeMask ? _GEN_1068 : _GEN_3116; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3629 = 4'h1 == io_writeMask ? _GEN_1069 : _GEN_3117; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3630 = 4'h1 == io_writeMask ? _GEN_1070 : _GEN_3118; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3631 = 4'h1 == io_writeMask ? _GEN_1071 : _GEN_3119; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3632 = 4'h1 == io_writeMask ? _GEN_1072 : _GEN_3120; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3633 = 4'h1 == io_writeMask ? _GEN_1073 : _GEN_3121; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3634 = 4'h1 == io_writeMask ? _GEN_1074 : _GEN_3122; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3635 = 4'h1 == io_writeMask ? _GEN_1075 : _GEN_3123; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3636 = 4'h1 == io_writeMask ? _GEN_1076 : _GEN_3124; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3637 = 4'h1 == io_writeMask ? _GEN_1077 : _GEN_3125; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3638 = 4'h1 == io_writeMask ? _GEN_1078 : _GEN_3126; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3639 = 4'h1 == io_writeMask ? _GEN_1079 : _GEN_3127; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3640 = 4'h1 == io_writeMask ? _GEN_1080 : _GEN_3128; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3641 = 4'h1 == io_writeMask ? _GEN_1081 : _GEN_3129; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3642 = 4'h1 == io_writeMask ? _GEN_1082 : _GEN_3130; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3643 = 4'h1 == io_writeMask ? _GEN_1083 : _GEN_3131; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3644 = 4'h1 == io_writeMask ? _GEN_1084 : _GEN_3132; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3645 = 4'h1 == io_writeMask ? _GEN_1085 : _GEN_3133; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3646 = 4'h1 == io_writeMask ? _GEN_1086 : _GEN_3134; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3647 = 4'h1 == io_writeMask ? _GEN_1087 : _GEN_3135; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3648 = 4'h1 == io_writeMask ? _GEN_1088 : _GEN_3136; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3649 = 4'h1 == io_writeMask ? _GEN_1089 : _GEN_3137; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3650 = 4'h1 == io_writeMask ? _GEN_1090 : _GEN_3138; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3651 = 4'h1 == io_writeMask ? _GEN_1091 : _GEN_3139; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3652 = 4'h1 == io_writeMask ? _GEN_1092 : _GEN_3140; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3653 = 4'h1 == io_writeMask ? _GEN_1093 : _GEN_3141; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3654 = 4'h1 == io_writeMask ? _GEN_1094 : _GEN_3142; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3655 = 4'h1 == io_writeMask ? _GEN_1095 : _GEN_3143; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3656 = 4'h1 == io_writeMask ? _GEN_1096 : _GEN_3144; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3657 = 4'h1 == io_writeMask ? _GEN_1097 : _GEN_3145; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3658 = 4'h1 == io_writeMask ? _GEN_1098 : _GEN_3146; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3659 = 4'h1 == io_writeMask ? _GEN_1099 : _GEN_3147; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3660 = 4'h1 == io_writeMask ? _GEN_1100 : _GEN_3148; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3661 = 4'h1 == io_writeMask ? _GEN_1101 : _GEN_3149; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3662 = 4'h1 == io_writeMask ? _GEN_1102 : _GEN_3150; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3663 = 4'h1 == io_writeMask ? _GEN_1103 : _GEN_3151; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3664 = 4'h1 == io_writeMask ? _GEN_1104 : _GEN_3152; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3665 = 4'h1 == io_writeMask ? _GEN_1105 : _GEN_3153; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3666 = 4'h1 == io_writeMask ? _GEN_1106 : _GEN_3154; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3667 = 4'h1 == io_writeMask ? _GEN_1107 : _GEN_3155; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3668 = 4'h1 == io_writeMask ? _GEN_1108 : _GEN_3156; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3669 = 4'h1 == io_writeMask ? _GEN_1109 : _GEN_3157; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3670 = 4'h1 == io_writeMask ? _GEN_1110 : _GEN_3158; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3671 = 4'h1 == io_writeMask ? _GEN_1111 : _GEN_3159; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3672 = 4'h1 == io_writeMask ? _GEN_1112 : _GEN_3160; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3673 = 4'h1 == io_writeMask ? _GEN_1113 : _GEN_3161; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3674 = 4'h1 == io_writeMask ? _GEN_1114 : _GEN_3162; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3675 = 4'h1 == io_writeMask ? _GEN_1115 : _GEN_3163; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3676 = 4'h1 == io_writeMask ? _GEN_1116 : _GEN_3164; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3677 = 4'h1 == io_writeMask ? _GEN_1117 : _GEN_3165; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3678 = 4'h1 == io_writeMask ? _GEN_1118 : _GEN_3166; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3679 = 4'h1 == io_writeMask ? _GEN_1119 : _GEN_3167; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3680 = 4'h1 == io_writeMask ? _GEN_1120 : _GEN_3168; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3681 = 4'h1 == io_writeMask ? _GEN_1121 : _GEN_3169; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3682 = 4'h1 == io_writeMask ? _GEN_1122 : _GEN_3170; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3683 = 4'h1 == io_writeMask ? _GEN_1123 : _GEN_3171; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3684 = 4'h1 == io_writeMask ? _GEN_1124 : _GEN_3172; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3685 = 4'h1 == io_writeMask ? _GEN_1125 : _GEN_3173; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3686 = 4'h1 == io_writeMask ? _GEN_1126 : _GEN_3174; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3687 = 4'h1 == io_writeMask ? _GEN_1127 : _GEN_3175; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3688 = 4'h1 == io_writeMask ? _GEN_1128 : _GEN_3176; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3689 = 4'h1 == io_writeMask ? _GEN_1129 : _GEN_3177; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3690 = 4'h1 == io_writeMask ? _GEN_1130 : _GEN_3178; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3691 = 4'h1 == io_writeMask ? _GEN_1131 : _GEN_3179; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3692 = 4'h1 == io_writeMask ? _GEN_1132 : _GEN_3180; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3693 = 4'h1 == io_writeMask ? _GEN_1133 : _GEN_3181; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3694 = 4'h1 == io_writeMask ? _GEN_1134 : _GEN_3182; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3695 = 4'h1 == io_writeMask ? _GEN_1135 : _GEN_3183; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3696 = 4'h1 == io_writeMask ? _GEN_1136 : _GEN_3184; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3697 = 4'h1 == io_writeMask ? _GEN_1137 : _GEN_3185; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3698 = 4'h1 == io_writeMask ? _GEN_1138 : _GEN_3186; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3699 = 4'h1 == io_writeMask ? _GEN_1139 : _GEN_3187; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3700 = 4'h1 == io_writeMask ? _GEN_1140 : _GEN_3188; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3701 = 4'h1 == io_writeMask ? _GEN_1141 : _GEN_3189; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3702 = 4'h1 == io_writeMask ? _GEN_1142 : _GEN_3190; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3703 = 4'h1 == io_writeMask ? _GEN_1143 : _GEN_3191; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3704 = 4'h1 == io_writeMask ? _GEN_1144 : _GEN_3192; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3705 = 4'h1 == io_writeMask ? _GEN_1145 : _GEN_3193; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3706 = 4'h1 == io_writeMask ? _GEN_1146 : _GEN_3194; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3707 = 4'h1 == io_writeMask ? _GEN_1147 : _GEN_3195; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3708 = 4'h1 == io_writeMask ? _GEN_1148 : _GEN_3196; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3709 = 4'h1 == io_writeMask ? _GEN_1149 : _GEN_3197; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3710 = 4'h1 == io_writeMask ? _GEN_1150 : _GEN_3198; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3711 = 4'h1 == io_writeMask ? _GEN_1151 : _GEN_3199; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3712 = 4'h1 == io_writeMask ? _GEN_1152 : _GEN_3200; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3713 = 4'h1 == io_writeMask ? _GEN_1153 : _GEN_3201; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3714 = 4'h1 == io_writeMask ? _GEN_1154 : _GEN_3202; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3715 = 4'h1 == io_writeMask ? _GEN_1155 : _GEN_3203; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3716 = 4'h1 == io_writeMask ? _GEN_1156 : _GEN_3204; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3717 = 4'h1 == io_writeMask ? _GEN_1157 : _GEN_3205; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3718 = 4'h1 == io_writeMask ? _GEN_1158 : _GEN_3206; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3719 = 4'h1 == io_writeMask ? _GEN_1159 : _GEN_3207; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3720 = 4'h1 == io_writeMask ? _GEN_1160 : _GEN_3208; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3721 = 4'h1 == io_writeMask ? _GEN_1161 : _GEN_3209; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3722 = 4'h1 == io_writeMask ? _GEN_1162 : _GEN_3210; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3723 = 4'h1 == io_writeMask ? _GEN_1163 : _GEN_3211; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3724 = 4'h1 == io_writeMask ? _GEN_1164 : _GEN_3212; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3725 = 4'h1 == io_writeMask ? _GEN_1165 : _GEN_3213; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3726 = 4'h1 == io_writeMask ? _GEN_1166 : _GEN_3214; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3727 = 4'h1 == io_writeMask ? _GEN_1167 : _GEN_3215; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3728 = 4'h1 == io_writeMask ? _GEN_1168 : _GEN_3216; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3729 = 4'h1 == io_writeMask ? _GEN_1169 : _GEN_3217; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3730 = 4'h1 == io_writeMask ? _GEN_1170 : _GEN_3218; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3731 = 4'h1 == io_writeMask ? _GEN_1171 : _GEN_3219; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3732 = 4'h1 == io_writeMask ? _GEN_1172 : _GEN_3220; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3733 = 4'h1 == io_writeMask ? _GEN_1173 : _GEN_3221; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3734 = 4'h1 == io_writeMask ? _GEN_1174 : _GEN_3222; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3735 = 4'h1 == io_writeMask ? _GEN_1175 : _GEN_3223; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3736 = 4'h1 == io_writeMask ? _GEN_1176 : _GEN_3224; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3737 = 4'h1 == io_writeMask ? _GEN_1177 : _GEN_3225; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3738 = 4'h1 == io_writeMask ? _GEN_1178 : _GEN_3226; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3739 = 4'h1 == io_writeMask ? _GEN_1179 : _GEN_3227; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3740 = 4'h1 == io_writeMask ? _GEN_1180 : _GEN_3228; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3741 = 4'h1 == io_writeMask ? _GEN_1181 : _GEN_3229; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3742 = 4'h1 == io_writeMask ? _GEN_1182 : _GEN_3230; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3743 = 4'h1 == io_writeMask ? _GEN_1183 : _GEN_3231; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3744 = 4'h1 == io_writeMask ? _GEN_1184 : _GEN_3232; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3745 = 4'h1 == io_writeMask ? _GEN_1185 : _GEN_3233; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3746 = 4'h1 == io_writeMask ? _GEN_1186 : _GEN_3234; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3747 = 4'h1 == io_writeMask ? _GEN_1187 : _GEN_3235; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3748 = 4'h1 == io_writeMask ? _GEN_1188 : _GEN_3236; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3749 = 4'h1 == io_writeMask ? _GEN_1189 : _GEN_3237; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3750 = 4'h1 == io_writeMask ? _GEN_1190 : _GEN_3238; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3751 = 4'h1 == io_writeMask ? _GEN_1191 : _GEN_3239; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3752 = 4'h1 == io_writeMask ? _GEN_1192 : _GEN_3240; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3753 = 4'h1 == io_writeMask ? _GEN_1193 : _GEN_3241; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3754 = 4'h1 == io_writeMask ? _GEN_1194 : _GEN_3242; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3755 = 4'h1 == io_writeMask ? _GEN_1195 : _GEN_3243; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3756 = 4'h1 == io_writeMask ? _GEN_1196 : _GEN_3244; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3757 = 4'h1 == io_writeMask ? _GEN_1197 : _GEN_3245; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3758 = 4'h1 == io_writeMask ? _GEN_1198 : _GEN_3246; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3759 = 4'h1 == io_writeMask ? _GEN_1199 : _GEN_3247; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3760 = 4'h1 == io_writeMask ? _GEN_1200 : _GEN_3248; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3761 = 4'h1 == io_writeMask ? _GEN_1201 : _GEN_3249; // @[Cache.scala 133:31]
  wire [31:0] _GEN_3762 = 4'h1 == io_writeMask ? _GEN_1202 : _GEN_3250; // @[Cache.scala 133:31]
  wire  _GEN_3763 = _GEN_9837 | dirty_0_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3764 = _GEN_9865 | dirty_0_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3765 = _GEN_9897 | dirty_0_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3766 = _GEN_9929 | dirty_0_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3767 = _GEN_9961 | dirty_0_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3768 = _GEN_9993 | dirty_0_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3769 = _GEN_10025 | dirty_0_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3770 = _GEN_10057 | dirty_0_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3771 = _GEN_10089 | dirty_1_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3772 = _GEN_10121 | dirty_1_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3773 = _GEN_10153 | dirty_1_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3774 = _GEN_10185 | dirty_1_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3775 = _GEN_10217 | dirty_1_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3776 = _GEN_10249 | dirty_1_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3777 = _GEN_10281 | dirty_1_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3778 = _GEN_10313 | dirty_1_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3779 = _GEN_10345 | dirty_2_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3780 = _GEN_10377 | dirty_2_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3781 = _GEN_10409 | dirty_2_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3782 = _GEN_10441 | dirty_2_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3783 = _GEN_10473 | dirty_2_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3784 = _GEN_10505 | dirty_2_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3785 = _GEN_10537 | dirty_2_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3786 = _GEN_10569 | dirty_2_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3787 = _GEN_10601 | dirty_3_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3788 = _GEN_10633 | dirty_3_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3789 = _GEN_10665 | dirty_3_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3790 = _GEN_10697 | dirty_3_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3791 = _GEN_10729 | dirty_3_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3792 = _GEN_10761 | dirty_3_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3793 = _GEN_10793 | dirty_3_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3794 = _GEN_10825 | dirty_3_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3795 = _GEN_10857 | dirty_4_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3796 = _GEN_10889 | dirty_4_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3797 = _GEN_10921 | dirty_4_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3798 = _GEN_10953 | dirty_4_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3799 = _GEN_10985 | dirty_4_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3800 = _GEN_11017 | dirty_4_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3801 = _GEN_11049 | dirty_4_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3802 = _GEN_11081 | dirty_4_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3803 = _GEN_11113 | dirty_5_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3804 = _GEN_11145 | dirty_5_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3805 = _GEN_11177 | dirty_5_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3806 = _GEN_11209 | dirty_5_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3807 = _GEN_11241 | dirty_5_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3808 = _GEN_11273 | dirty_5_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3809 = _GEN_11305 | dirty_5_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3810 = _GEN_11337 | dirty_5_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3811 = _GEN_11369 | dirty_6_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3812 = _GEN_11401 | dirty_6_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3813 = _GEN_11433 | dirty_6_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3814 = _GEN_11465 | dirty_6_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3815 = _GEN_11497 | dirty_6_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3816 = _GEN_11529 | dirty_6_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3817 = _GEN_11561 | dirty_6_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3818 = _GEN_11593 | dirty_6_7; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3819 = _GEN_11625 | dirty_7_0; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3820 = _GEN_11657 | dirty_7_1; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3821 = _GEN_11689 | dirty_7_2; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3822 = _GEN_11721 | dirty_7_3; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3823 = _GEN_11753 | dirty_7_4; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3824 = _GEN_11785 | dirty_7_5; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3825 = _GEN_11817 | dirty_7_6; // @[Cache.scala 144:{36,36} 58:22]
  wire  _GEN_3826 = _GEN_11849 | dirty_7_7; // @[Cache.scala 144:{36,36} 58:22]
  wire [31:0] _GEN_3827 = io_w_req ? _GEN_3251 : CacheMem_0_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3828 = io_w_req ? _GEN_3252 : CacheMem_0_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3829 = io_w_req ? _GEN_3253 : CacheMem_0_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3830 = io_w_req ? _GEN_3254 : CacheMem_0_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3831 = io_w_req ? _GEN_3255 : CacheMem_0_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3832 = io_w_req ? _GEN_3256 : CacheMem_0_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3833 = io_w_req ? _GEN_3257 : CacheMem_0_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3834 = io_w_req ? _GEN_3258 : CacheMem_0_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3835 = io_w_req ? _GEN_3259 : CacheMem_0_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3836 = io_w_req ? _GEN_3260 : CacheMem_0_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3837 = io_w_req ? _GEN_3261 : CacheMem_0_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3838 = io_w_req ? _GEN_3262 : CacheMem_0_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3839 = io_w_req ? _GEN_3263 : CacheMem_0_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3840 = io_w_req ? _GEN_3264 : CacheMem_0_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3841 = io_w_req ? _GEN_3265 : CacheMem_0_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3842 = io_w_req ? _GEN_3266 : CacheMem_0_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3843 = io_w_req ? _GEN_3267 : CacheMem_0_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3844 = io_w_req ? _GEN_3268 : CacheMem_0_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3845 = io_w_req ? _GEN_3269 : CacheMem_0_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3846 = io_w_req ? _GEN_3270 : CacheMem_0_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3847 = io_w_req ? _GEN_3271 : CacheMem_0_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3848 = io_w_req ? _GEN_3272 : CacheMem_0_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3849 = io_w_req ? _GEN_3273 : CacheMem_0_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3850 = io_w_req ? _GEN_3274 : CacheMem_0_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3851 = io_w_req ? _GEN_3275 : CacheMem_0_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3852 = io_w_req ? _GEN_3276 : CacheMem_0_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3853 = io_w_req ? _GEN_3277 : CacheMem_0_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3854 = io_w_req ? _GEN_3278 : CacheMem_0_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3855 = io_w_req ? _GEN_3279 : CacheMem_0_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3856 = io_w_req ? _GEN_3280 : CacheMem_0_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3857 = io_w_req ? _GEN_3281 : CacheMem_0_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3858 = io_w_req ? _GEN_3282 : CacheMem_0_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3859 = io_w_req ? _GEN_3283 : CacheMem_0_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3860 = io_w_req ? _GEN_3284 : CacheMem_0_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3861 = io_w_req ? _GEN_3285 : CacheMem_0_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3862 = io_w_req ? _GEN_3286 : CacheMem_0_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3863 = io_w_req ? _GEN_3287 : CacheMem_0_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3864 = io_w_req ? _GEN_3288 : CacheMem_0_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3865 = io_w_req ? _GEN_3289 : CacheMem_0_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3866 = io_w_req ? _GEN_3290 : CacheMem_0_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3867 = io_w_req ? _GEN_3291 : CacheMem_0_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3868 = io_w_req ? _GEN_3292 : CacheMem_0_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3869 = io_w_req ? _GEN_3293 : CacheMem_0_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3870 = io_w_req ? _GEN_3294 : CacheMem_0_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3871 = io_w_req ? _GEN_3295 : CacheMem_0_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3872 = io_w_req ? _GEN_3296 : CacheMem_0_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3873 = io_w_req ? _GEN_3297 : CacheMem_0_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3874 = io_w_req ? _GEN_3298 : CacheMem_0_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3875 = io_w_req ? _GEN_3299 : CacheMem_0_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3876 = io_w_req ? _GEN_3300 : CacheMem_0_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3877 = io_w_req ? _GEN_3301 : CacheMem_0_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3878 = io_w_req ? _GEN_3302 : CacheMem_0_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3879 = io_w_req ? _GEN_3303 : CacheMem_0_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3880 = io_w_req ? _GEN_3304 : CacheMem_0_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3881 = io_w_req ? _GEN_3305 : CacheMem_0_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3882 = io_w_req ? _GEN_3306 : CacheMem_0_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3883 = io_w_req ? _GEN_3307 : CacheMem_0_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3884 = io_w_req ? _GEN_3308 : CacheMem_0_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3885 = io_w_req ? _GEN_3309 : CacheMem_0_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3886 = io_w_req ? _GEN_3310 : CacheMem_0_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3887 = io_w_req ? _GEN_3311 : CacheMem_0_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3888 = io_w_req ? _GEN_3312 : CacheMem_0_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3889 = io_w_req ? _GEN_3313 : CacheMem_0_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3890 = io_w_req ? _GEN_3314 : CacheMem_0_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3891 = io_w_req ? _GEN_3315 : CacheMem_1_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3892 = io_w_req ? _GEN_3316 : CacheMem_1_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3893 = io_w_req ? _GEN_3317 : CacheMem_1_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3894 = io_w_req ? _GEN_3318 : CacheMem_1_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3895 = io_w_req ? _GEN_3319 : CacheMem_1_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3896 = io_w_req ? _GEN_3320 : CacheMem_1_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3897 = io_w_req ? _GEN_3321 : CacheMem_1_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3898 = io_w_req ? _GEN_3322 : CacheMem_1_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3899 = io_w_req ? _GEN_3323 : CacheMem_1_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3900 = io_w_req ? _GEN_3324 : CacheMem_1_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3901 = io_w_req ? _GEN_3325 : CacheMem_1_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3902 = io_w_req ? _GEN_3326 : CacheMem_1_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3903 = io_w_req ? _GEN_3327 : CacheMem_1_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3904 = io_w_req ? _GEN_3328 : CacheMem_1_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3905 = io_w_req ? _GEN_3329 : CacheMem_1_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3906 = io_w_req ? _GEN_3330 : CacheMem_1_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3907 = io_w_req ? _GEN_3331 : CacheMem_1_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3908 = io_w_req ? _GEN_3332 : CacheMem_1_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3909 = io_w_req ? _GEN_3333 : CacheMem_1_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3910 = io_w_req ? _GEN_3334 : CacheMem_1_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3911 = io_w_req ? _GEN_3335 : CacheMem_1_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3912 = io_w_req ? _GEN_3336 : CacheMem_1_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3913 = io_w_req ? _GEN_3337 : CacheMem_1_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3914 = io_w_req ? _GEN_3338 : CacheMem_1_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3915 = io_w_req ? _GEN_3339 : CacheMem_1_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3916 = io_w_req ? _GEN_3340 : CacheMem_1_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3917 = io_w_req ? _GEN_3341 : CacheMem_1_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3918 = io_w_req ? _GEN_3342 : CacheMem_1_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3919 = io_w_req ? _GEN_3343 : CacheMem_1_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3920 = io_w_req ? _GEN_3344 : CacheMem_1_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3921 = io_w_req ? _GEN_3345 : CacheMem_1_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3922 = io_w_req ? _GEN_3346 : CacheMem_1_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3923 = io_w_req ? _GEN_3347 : CacheMem_1_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3924 = io_w_req ? _GEN_3348 : CacheMem_1_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3925 = io_w_req ? _GEN_3349 : CacheMem_1_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3926 = io_w_req ? _GEN_3350 : CacheMem_1_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3927 = io_w_req ? _GEN_3351 : CacheMem_1_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3928 = io_w_req ? _GEN_3352 : CacheMem_1_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3929 = io_w_req ? _GEN_3353 : CacheMem_1_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3930 = io_w_req ? _GEN_3354 : CacheMem_1_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3931 = io_w_req ? _GEN_3355 : CacheMem_1_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3932 = io_w_req ? _GEN_3356 : CacheMem_1_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3933 = io_w_req ? _GEN_3357 : CacheMem_1_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3934 = io_w_req ? _GEN_3358 : CacheMem_1_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3935 = io_w_req ? _GEN_3359 : CacheMem_1_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3936 = io_w_req ? _GEN_3360 : CacheMem_1_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3937 = io_w_req ? _GEN_3361 : CacheMem_1_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3938 = io_w_req ? _GEN_3362 : CacheMem_1_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3939 = io_w_req ? _GEN_3363 : CacheMem_1_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3940 = io_w_req ? _GEN_3364 : CacheMem_1_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3941 = io_w_req ? _GEN_3365 : CacheMem_1_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3942 = io_w_req ? _GEN_3366 : CacheMem_1_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3943 = io_w_req ? _GEN_3367 : CacheMem_1_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3944 = io_w_req ? _GEN_3368 : CacheMem_1_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3945 = io_w_req ? _GEN_3369 : CacheMem_1_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3946 = io_w_req ? _GEN_3370 : CacheMem_1_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3947 = io_w_req ? _GEN_3371 : CacheMem_1_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3948 = io_w_req ? _GEN_3372 : CacheMem_1_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3949 = io_w_req ? _GEN_3373 : CacheMem_1_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3950 = io_w_req ? _GEN_3374 : CacheMem_1_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3951 = io_w_req ? _GEN_3375 : CacheMem_1_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3952 = io_w_req ? _GEN_3376 : CacheMem_1_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3953 = io_w_req ? _GEN_3377 : CacheMem_1_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3954 = io_w_req ? _GEN_3378 : CacheMem_1_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3955 = io_w_req ? _GEN_3379 : CacheMem_2_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3956 = io_w_req ? _GEN_3380 : CacheMem_2_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3957 = io_w_req ? _GEN_3381 : CacheMem_2_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3958 = io_w_req ? _GEN_3382 : CacheMem_2_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3959 = io_w_req ? _GEN_3383 : CacheMem_2_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3960 = io_w_req ? _GEN_3384 : CacheMem_2_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3961 = io_w_req ? _GEN_3385 : CacheMem_2_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3962 = io_w_req ? _GEN_3386 : CacheMem_2_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3963 = io_w_req ? _GEN_3387 : CacheMem_2_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3964 = io_w_req ? _GEN_3388 : CacheMem_2_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3965 = io_w_req ? _GEN_3389 : CacheMem_2_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3966 = io_w_req ? _GEN_3390 : CacheMem_2_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3967 = io_w_req ? _GEN_3391 : CacheMem_2_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3968 = io_w_req ? _GEN_3392 : CacheMem_2_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3969 = io_w_req ? _GEN_3393 : CacheMem_2_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3970 = io_w_req ? _GEN_3394 : CacheMem_2_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3971 = io_w_req ? _GEN_3395 : CacheMem_2_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3972 = io_w_req ? _GEN_3396 : CacheMem_2_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3973 = io_w_req ? _GEN_3397 : CacheMem_2_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3974 = io_w_req ? _GEN_3398 : CacheMem_2_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3975 = io_w_req ? _GEN_3399 : CacheMem_2_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3976 = io_w_req ? _GEN_3400 : CacheMem_2_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3977 = io_w_req ? _GEN_3401 : CacheMem_2_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3978 = io_w_req ? _GEN_3402 : CacheMem_2_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3979 = io_w_req ? _GEN_3403 : CacheMem_2_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3980 = io_w_req ? _GEN_3404 : CacheMem_2_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3981 = io_w_req ? _GEN_3405 : CacheMem_2_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3982 = io_w_req ? _GEN_3406 : CacheMem_2_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3983 = io_w_req ? _GEN_3407 : CacheMem_2_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3984 = io_w_req ? _GEN_3408 : CacheMem_2_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3985 = io_w_req ? _GEN_3409 : CacheMem_2_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3986 = io_w_req ? _GEN_3410 : CacheMem_2_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3987 = io_w_req ? _GEN_3411 : CacheMem_2_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3988 = io_w_req ? _GEN_3412 : CacheMem_2_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3989 = io_w_req ? _GEN_3413 : CacheMem_2_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3990 = io_w_req ? _GEN_3414 : CacheMem_2_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3991 = io_w_req ? _GEN_3415 : CacheMem_2_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3992 = io_w_req ? _GEN_3416 : CacheMem_2_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3993 = io_w_req ? _GEN_3417 : CacheMem_2_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3994 = io_w_req ? _GEN_3418 : CacheMem_2_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3995 = io_w_req ? _GEN_3419 : CacheMem_2_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3996 = io_w_req ? _GEN_3420 : CacheMem_2_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3997 = io_w_req ? _GEN_3421 : CacheMem_2_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3998 = io_w_req ? _GEN_3422 : CacheMem_2_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_3999 = io_w_req ? _GEN_3423 : CacheMem_2_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4000 = io_w_req ? _GEN_3424 : CacheMem_2_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4001 = io_w_req ? _GEN_3425 : CacheMem_2_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4002 = io_w_req ? _GEN_3426 : CacheMem_2_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4003 = io_w_req ? _GEN_3427 : CacheMem_2_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4004 = io_w_req ? _GEN_3428 : CacheMem_2_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4005 = io_w_req ? _GEN_3429 : CacheMem_2_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4006 = io_w_req ? _GEN_3430 : CacheMem_2_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4007 = io_w_req ? _GEN_3431 : CacheMem_2_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4008 = io_w_req ? _GEN_3432 : CacheMem_2_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4009 = io_w_req ? _GEN_3433 : CacheMem_2_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4010 = io_w_req ? _GEN_3434 : CacheMem_2_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4011 = io_w_req ? _GEN_3435 : CacheMem_2_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4012 = io_w_req ? _GEN_3436 : CacheMem_2_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4013 = io_w_req ? _GEN_3437 : CacheMem_2_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4014 = io_w_req ? _GEN_3438 : CacheMem_2_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4015 = io_w_req ? _GEN_3439 : CacheMem_2_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4016 = io_w_req ? _GEN_3440 : CacheMem_2_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4017 = io_w_req ? _GEN_3441 : CacheMem_2_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4018 = io_w_req ? _GEN_3442 : CacheMem_2_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4019 = io_w_req ? _GEN_3443 : CacheMem_3_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4020 = io_w_req ? _GEN_3444 : CacheMem_3_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4021 = io_w_req ? _GEN_3445 : CacheMem_3_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4022 = io_w_req ? _GEN_3446 : CacheMem_3_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4023 = io_w_req ? _GEN_3447 : CacheMem_3_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4024 = io_w_req ? _GEN_3448 : CacheMem_3_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4025 = io_w_req ? _GEN_3449 : CacheMem_3_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4026 = io_w_req ? _GEN_3450 : CacheMem_3_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4027 = io_w_req ? _GEN_3451 : CacheMem_3_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4028 = io_w_req ? _GEN_3452 : CacheMem_3_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4029 = io_w_req ? _GEN_3453 : CacheMem_3_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4030 = io_w_req ? _GEN_3454 : CacheMem_3_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4031 = io_w_req ? _GEN_3455 : CacheMem_3_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4032 = io_w_req ? _GEN_3456 : CacheMem_3_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4033 = io_w_req ? _GEN_3457 : CacheMem_3_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4034 = io_w_req ? _GEN_3458 : CacheMem_3_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4035 = io_w_req ? _GEN_3459 : CacheMem_3_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4036 = io_w_req ? _GEN_3460 : CacheMem_3_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4037 = io_w_req ? _GEN_3461 : CacheMem_3_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4038 = io_w_req ? _GEN_3462 : CacheMem_3_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4039 = io_w_req ? _GEN_3463 : CacheMem_3_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4040 = io_w_req ? _GEN_3464 : CacheMem_3_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4041 = io_w_req ? _GEN_3465 : CacheMem_3_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4042 = io_w_req ? _GEN_3466 : CacheMem_3_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4043 = io_w_req ? _GEN_3467 : CacheMem_3_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4044 = io_w_req ? _GEN_3468 : CacheMem_3_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4045 = io_w_req ? _GEN_3469 : CacheMem_3_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4046 = io_w_req ? _GEN_3470 : CacheMem_3_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4047 = io_w_req ? _GEN_3471 : CacheMem_3_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4048 = io_w_req ? _GEN_3472 : CacheMem_3_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4049 = io_w_req ? _GEN_3473 : CacheMem_3_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4050 = io_w_req ? _GEN_3474 : CacheMem_3_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4051 = io_w_req ? _GEN_3475 : CacheMem_3_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4052 = io_w_req ? _GEN_3476 : CacheMem_3_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4053 = io_w_req ? _GEN_3477 : CacheMem_3_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4054 = io_w_req ? _GEN_3478 : CacheMem_3_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4055 = io_w_req ? _GEN_3479 : CacheMem_3_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4056 = io_w_req ? _GEN_3480 : CacheMem_3_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4057 = io_w_req ? _GEN_3481 : CacheMem_3_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4058 = io_w_req ? _GEN_3482 : CacheMem_3_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4059 = io_w_req ? _GEN_3483 : CacheMem_3_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4060 = io_w_req ? _GEN_3484 : CacheMem_3_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4061 = io_w_req ? _GEN_3485 : CacheMem_3_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4062 = io_w_req ? _GEN_3486 : CacheMem_3_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4063 = io_w_req ? _GEN_3487 : CacheMem_3_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4064 = io_w_req ? _GEN_3488 : CacheMem_3_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4065 = io_w_req ? _GEN_3489 : CacheMem_3_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4066 = io_w_req ? _GEN_3490 : CacheMem_3_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4067 = io_w_req ? _GEN_3491 : CacheMem_3_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4068 = io_w_req ? _GEN_3492 : CacheMem_3_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4069 = io_w_req ? _GEN_3493 : CacheMem_3_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4070 = io_w_req ? _GEN_3494 : CacheMem_3_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4071 = io_w_req ? _GEN_3495 : CacheMem_3_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4072 = io_w_req ? _GEN_3496 : CacheMem_3_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4073 = io_w_req ? _GEN_3497 : CacheMem_3_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4074 = io_w_req ? _GEN_3498 : CacheMem_3_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4075 = io_w_req ? _GEN_3499 : CacheMem_3_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4076 = io_w_req ? _GEN_3500 : CacheMem_3_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4077 = io_w_req ? _GEN_3501 : CacheMem_3_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4078 = io_w_req ? _GEN_3502 : CacheMem_3_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4079 = io_w_req ? _GEN_3503 : CacheMem_3_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4080 = io_w_req ? _GEN_3504 : CacheMem_3_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4081 = io_w_req ? _GEN_3505 : CacheMem_3_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4082 = io_w_req ? _GEN_3506 : CacheMem_3_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4083 = io_w_req ? _GEN_3507 : CacheMem_4_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4084 = io_w_req ? _GEN_3508 : CacheMem_4_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4085 = io_w_req ? _GEN_3509 : CacheMem_4_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4086 = io_w_req ? _GEN_3510 : CacheMem_4_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4087 = io_w_req ? _GEN_3511 : CacheMem_4_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4088 = io_w_req ? _GEN_3512 : CacheMem_4_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4089 = io_w_req ? _GEN_3513 : CacheMem_4_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4090 = io_w_req ? _GEN_3514 : CacheMem_4_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4091 = io_w_req ? _GEN_3515 : CacheMem_4_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4092 = io_w_req ? _GEN_3516 : CacheMem_4_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4093 = io_w_req ? _GEN_3517 : CacheMem_4_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4094 = io_w_req ? _GEN_3518 : CacheMem_4_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4095 = io_w_req ? _GEN_3519 : CacheMem_4_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4096 = io_w_req ? _GEN_3520 : CacheMem_4_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4097 = io_w_req ? _GEN_3521 : CacheMem_4_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4098 = io_w_req ? _GEN_3522 : CacheMem_4_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4099 = io_w_req ? _GEN_3523 : CacheMem_4_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4100 = io_w_req ? _GEN_3524 : CacheMem_4_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4101 = io_w_req ? _GEN_3525 : CacheMem_4_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4102 = io_w_req ? _GEN_3526 : CacheMem_4_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4103 = io_w_req ? _GEN_3527 : CacheMem_4_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4104 = io_w_req ? _GEN_3528 : CacheMem_4_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4105 = io_w_req ? _GEN_3529 : CacheMem_4_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4106 = io_w_req ? _GEN_3530 : CacheMem_4_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4107 = io_w_req ? _GEN_3531 : CacheMem_4_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4108 = io_w_req ? _GEN_3532 : CacheMem_4_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4109 = io_w_req ? _GEN_3533 : CacheMem_4_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4110 = io_w_req ? _GEN_3534 : CacheMem_4_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4111 = io_w_req ? _GEN_3535 : CacheMem_4_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4112 = io_w_req ? _GEN_3536 : CacheMem_4_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4113 = io_w_req ? _GEN_3537 : CacheMem_4_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4114 = io_w_req ? _GEN_3538 : CacheMem_4_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4115 = io_w_req ? _GEN_3539 : CacheMem_4_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4116 = io_w_req ? _GEN_3540 : CacheMem_4_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4117 = io_w_req ? _GEN_3541 : CacheMem_4_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4118 = io_w_req ? _GEN_3542 : CacheMem_4_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4119 = io_w_req ? _GEN_3543 : CacheMem_4_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4120 = io_w_req ? _GEN_3544 : CacheMem_4_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4121 = io_w_req ? _GEN_3545 : CacheMem_4_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4122 = io_w_req ? _GEN_3546 : CacheMem_4_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4123 = io_w_req ? _GEN_3547 : CacheMem_4_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4124 = io_w_req ? _GEN_3548 : CacheMem_4_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4125 = io_w_req ? _GEN_3549 : CacheMem_4_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4126 = io_w_req ? _GEN_3550 : CacheMem_4_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4127 = io_w_req ? _GEN_3551 : CacheMem_4_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4128 = io_w_req ? _GEN_3552 : CacheMem_4_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4129 = io_w_req ? _GEN_3553 : CacheMem_4_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4130 = io_w_req ? _GEN_3554 : CacheMem_4_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4131 = io_w_req ? _GEN_3555 : CacheMem_4_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4132 = io_w_req ? _GEN_3556 : CacheMem_4_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4133 = io_w_req ? _GEN_3557 : CacheMem_4_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4134 = io_w_req ? _GEN_3558 : CacheMem_4_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4135 = io_w_req ? _GEN_3559 : CacheMem_4_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4136 = io_w_req ? _GEN_3560 : CacheMem_4_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4137 = io_w_req ? _GEN_3561 : CacheMem_4_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4138 = io_w_req ? _GEN_3562 : CacheMem_4_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4139 = io_w_req ? _GEN_3563 : CacheMem_4_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4140 = io_w_req ? _GEN_3564 : CacheMem_4_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4141 = io_w_req ? _GEN_3565 : CacheMem_4_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4142 = io_w_req ? _GEN_3566 : CacheMem_4_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4143 = io_w_req ? _GEN_3567 : CacheMem_4_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4144 = io_w_req ? _GEN_3568 : CacheMem_4_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4145 = io_w_req ? _GEN_3569 : CacheMem_4_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4146 = io_w_req ? _GEN_3570 : CacheMem_4_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4147 = io_w_req ? _GEN_3571 : CacheMem_5_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4148 = io_w_req ? _GEN_3572 : CacheMem_5_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4149 = io_w_req ? _GEN_3573 : CacheMem_5_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4150 = io_w_req ? _GEN_3574 : CacheMem_5_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4151 = io_w_req ? _GEN_3575 : CacheMem_5_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4152 = io_w_req ? _GEN_3576 : CacheMem_5_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4153 = io_w_req ? _GEN_3577 : CacheMem_5_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4154 = io_w_req ? _GEN_3578 : CacheMem_5_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4155 = io_w_req ? _GEN_3579 : CacheMem_5_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4156 = io_w_req ? _GEN_3580 : CacheMem_5_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4157 = io_w_req ? _GEN_3581 : CacheMem_5_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4158 = io_w_req ? _GEN_3582 : CacheMem_5_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4159 = io_w_req ? _GEN_3583 : CacheMem_5_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4160 = io_w_req ? _GEN_3584 : CacheMem_5_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4161 = io_w_req ? _GEN_3585 : CacheMem_5_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4162 = io_w_req ? _GEN_3586 : CacheMem_5_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4163 = io_w_req ? _GEN_3587 : CacheMem_5_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4164 = io_w_req ? _GEN_3588 : CacheMem_5_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4165 = io_w_req ? _GEN_3589 : CacheMem_5_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4166 = io_w_req ? _GEN_3590 : CacheMem_5_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4167 = io_w_req ? _GEN_3591 : CacheMem_5_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4168 = io_w_req ? _GEN_3592 : CacheMem_5_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4169 = io_w_req ? _GEN_3593 : CacheMem_5_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4170 = io_w_req ? _GEN_3594 : CacheMem_5_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4171 = io_w_req ? _GEN_3595 : CacheMem_5_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4172 = io_w_req ? _GEN_3596 : CacheMem_5_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4173 = io_w_req ? _GEN_3597 : CacheMem_5_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4174 = io_w_req ? _GEN_3598 : CacheMem_5_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4175 = io_w_req ? _GEN_3599 : CacheMem_5_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4176 = io_w_req ? _GEN_3600 : CacheMem_5_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4177 = io_w_req ? _GEN_3601 : CacheMem_5_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4178 = io_w_req ? _GEN_3602 : CacheMem_5_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4179 = io_w_req ? _GEN_3603 : CacheMem_5_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4180 = io_w_req ? _GEN_3604 : CacheMem_5_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4181 = io_w_req ? _GEN_3605 : CacheMem_5_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4182 = io_w_req ? _GEN_3606 : CacheMem_5_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4183 = io_w_req ? _GEN_3607 : CacheMem_5_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4184 = io_w_req ? _GEN_3608 : CacheMem_5_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4185 = io_w_req ? _GEN_3609 : CacheMem_5_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4186 = io_w_req ? _GEN_3610 : CacheMem_5_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4187 = io_w_req ? _GEN_3611 : CacheMem_5_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4188 = io_w_req ? _GEN_3612 : CacheMem_5_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4189 = io_w_req ? _GEN_3613 : CacheMem_5_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4190 = io_w_req ? _GEN_3614 : CacheMem_5_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4191 = io_w_req ? _GEN_3615 : CacheMem_5_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4192 = io_w_req ? _GEN_3616 : CacheMem_5_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4193 = io_w_req ? _GEN_3617 : CacheMem_5_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4194 = io_w_req ? _GEN_3618 : CacheMem_5_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4195 = io_w_req ? _GEN_3619 : CacheMem_5_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4196 = io_w_req ? _GEN_3620 : CacheMem_5_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4197 = io_w_req ? _GEN_3621 : CacheMem_5_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4198 = io_w_req ? _GEN_3622 : CacheMem_5_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4199 = io_w_req ? _GEN_3623 : CacheMem_5_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4200 = io_w_req ? _GEN_3624 : CacheMem_5_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4201 = io_w_req ? _GEN_3625 : CacheMem_5_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4202 = io_w_req ? _GEN_3626 : CacheMem_5_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4203 = io_w_req ? _GEN_3627 : CacheMem_5_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4204 = io_w_req ? _GEN_3628 : CacheMem_5_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4205 = io_w_req ? _GEN_3629 : CacheMem_5_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4206 = io_w_req ? _GEN_3630 : CacheMem_5_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4207 = io_w_req ? _GEN_3631 : CacheMem_5_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4208 = io_w_req ? _GEN_3632 : CacheMem_5_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4209 = io_w_req ? _GEN_3633 : CacheMem_5_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4210 = io_w_req ? _GEN_3634 : CacheMem_5_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4211 = io_w_req ? _GEN_3635 : CacheMem_6_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4212 = io_w_req ? _GEN_3636 : CacheMem_6_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4213 = io_w_req ? _GEN_3637 : CacheMem_6_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4214 = io_w_req ? _GEN_3638 : CacheMem_6_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4215 = io_w_req ? _GEN_3639 : CacheMem_6_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4216 = io_w_req ? _GEN_3640 : CacheMem_6_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4217 = io_w_req ? _GEN_3641 : CacheMem_6_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4218 = io_w_req ? _GEN_3642 : CacheMem_6_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4219 = io_w_req ? _GEN_3643 : CacheMem_6_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4220 = io_w_req ? _GEN_3644 : CacheMem_6_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4221 = io_w_req ? _GEN_3645 : CacheMem_6_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4222 = io_w_req ? _GEN_3646 : CacheMem_6_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4223 = io_w_req ? _GEN_3647 : CacheMem_6_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4224 = io_w_req ? _GEN_3648 : CacheMem_6_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4225 = io_w_req ? _GEN_3649 : CacheMem_6_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4226 = io_w_req ? _GEN_3650 : CacheMem_6_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4227 = io_w_req ? _GEN_3651 : CacheMem_6_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4228 = io_w_req ? _GEN_3652 : CacheMem_6_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4229 = io_w_req ? _GEN_3653 : CacheMem_6_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4230 = io_w_req ? _GEN_3654 : CacheMem_6_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4231 = io_w_req ? _GEN_3655 : CacheMem_6_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4232 = io_w_req ? _GEN_3656 : CacheMem_6_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4233 = io_w_req ? _GEN_3657 : CacheMem_6_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4234 = io_w_req ? _GEN_3658 : CacheMem_6_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4235 = io_w_req ? _GEN_3659 : CacheMem_6_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4236 = io_w_req ? _GEN_3660 : CacheMem_6_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4237 = io_w_req ? _GEN_3661 : CacheMem_6_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4238 = io_w_req ? _GEN_3662 : CacheMem_6_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4239 = io_w_req ? _GEN_3663 : CacheMem_6_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4240 = io_w_req ? _GEN_3664 : CacheMem_6_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4241 = io_w_req ? _GEN_3665 : CacheMem_6_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4242 = io_w_req ? _GEN_3666 : CacheMem_6_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4243 = io_w_req ? _GEN_3667 : CacheMem_6_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4244 = io_w_req ? _GEN_3668 : CacheMem_6_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4245 = io_w_req ? _GEN_3669 : CacheMem_6_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4246 = io_w_req ? _GEN_3670 : CacheMem_6_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4247 = io_w_req ? _GEN_3671 : CacheMem_6_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4248 = io_w_req ? _GEN_3672 : CacheMem_6_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4249 = io_w_req ? _GEN_3673 : CacheMem_6_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4250 = io_w_req ? _GEN_3674 : CacheMem_6_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4251 = io_w_req ? _GEN_3675 : CacheMem_6_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4252 = io_w_req ? _GEN_3676 : CacheMem_6_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4253 = io_w_req ? _GEN_3677 : CacheMem_6_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4254 = io_w_req ? _GEN_3678 : CacheMem_6_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4255 = io_w_req ? _GEN_3679 : CacheMem_6_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4256 = io_w_req ? _GEN_3680 : CacheMem_6_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4257 = io_w_req ? _GEN_3681 : CacheMem_6_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4258 = io_w_req ? _GEN_3682 : CacheMem_6_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4259 = io_w_req ? _GEN_3683 : CacheMem_6_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4260 = io_w_req ? _GEN_3684 : CacheMem_6_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4261 = io_w_req ? _GEN_3685 : CacheMem_6_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4262 = io_w_req ? _GEN_3686 : CacheMem_6_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4263 = io_w_req ? _GEN_3687 : CacheMem_6_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4264 = io_w_req ? _GEN_3688 : CacheMem_6_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4265 = io_w_req ? _GEN_3689 : CacheMem_6_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4266 = io_w_req ? _GEN_3690 : CacheMem_6_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4267 = io_w_req ? _GEN_3691 : CacheMem_6_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4268 = io_w_req ? _GEN_3692 : CacheMem_6_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4269 = io_w_req ? _GEN_3693 : CacheMem_6_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4270 = io_w_req ? _GEN_3694 : CacheMem_6_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4271 = io_w_req ? _GEN_3695 : CacheMem_6_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4272 = io_w_req ? _GEN_3696 : CacheMem_6_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4273 = io_w_req ? _GEN_3697 : CacheMem_6_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4274 = io_w_req ? _GEN_3698 : CacheMem_6_7_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4275 = io_w_req ? _GEN_3699 : CacheMem_7_0_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4276 = io_w_req ? _GEN_3700 : CacheMem_7_0_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4277 = io_w_req ? _GEN_3701 : CacheMem_7_0_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4278 = io_w_req ? _GEN_3702 : CacheMem_7_0_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4279 = io_w_req ? _GEN_3703 : CacheMem_7_0_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4280 = io_w_req ? _GEN_3704 : CacheMem_7_0_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4281 = io_w_req ? _GEN_3705 : CacheMem_7_0_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4282 = io_w_req ? _GEN_3706 : CacheMem_7_0_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4283 = io_w_req ? _GEN_3707 : CacheMem_7_1_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4284 = io_w_req ? _GEN_3708 : CacheMem_7_1_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4285 = io_w_req ? _GEN_3709 : CacheMem_7_1_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4286 = io_w_req ? _GEN_3710 : CacheMem_7_1_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4287 = io_w_req ? _GEN_3711 : CacheMem_7_1_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4288 = io_w_req ? _GEN_3712 : CacheMem_7_1_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4289 = io_w_req ? _GEN_3713 : CacheMem_7_1_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4290 = io_w_req ? _GEN_3714 : CacheMem_7_1_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4291 = io_w_req ? _GEN_3715 : CacheMem_7_2_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4292 = io_w_req ? _GEN_3716 : CacheMem_7_2_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4293 = io_w_req ? _GEN_3717 : CacheMem_7_2_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4294 = io_w_req ? _GEN_3718 : CacheMem_7_2_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4295 = io_w_req ? _GEN_3719 : CacheMem_7_2_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4296 = io_w_req ? _GEN_3720 : CacheMem_7_2_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4297 = io_w_req ? _GEN_3721 : CacheMem_7_2_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4298 = io_w_req ? _GEN_3722 : CacheMem_7_2_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4299 = io_w_req ? _GEN_3723 : CacheMem_7_3_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4300 = io_w_req ? _GEN_3724 : CacheMem_7_3_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4301 = io_w_req ? _GEN_3725 : CacheMem_7_3_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4302 = io_w_req ? _GEN_3726 : CacheMem_7_3_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4303 = io_w_req ? _GEN_3727 : CacheMem_7_3_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4304 = io_w_req ? _GEN_3728 : CacheMem_7_3_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4305 = io_w_req ? _GEN_3729 : CacheMem_7_3_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4306 = io_w_req ? _GEN_3730 : CacheMem_7_3_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4307 = io_w_req ? _GEN_3731 : CacheMem_7_4_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4308 = io_w_req ? _GEN_3732 : CacheMem_7_4_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4309 = io_w_req ? _GEN_3733 : CacheMem_7_4_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4310 = io_w_req ? _GEN_3734 : CacheMem_7_4_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4311 = io_w_req ? _GEN_3735 : CacheMem_7_4_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4312 = io_w_req ? _GEN_3736 : CacheMem_7_4_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4313 = io_w_req ? _GEN_3737 : CacheMem_7_4_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4314 = io_w_req ? _GEN_3738 : CacheMem_7_4_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4315 = io_w_req ? _GEN_3739 : CacheMem_7_5_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4316 = io_w_req ? _GEN_3740 : CacheMem_7_5_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4317 = io_w_req ? _GEN_3741 : CacheMem_7_5_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4318 = io_w_req ? _GEN_3742 : CacheMem_7_5_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4319 = io_w_req ? _GEN_3743 : CacheMem_7_5_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4320 = io_w_req ? _GEN_3744 : CacheMem_7_5_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4321 = io_w_req ? _GEN_3745 : CacheMem_7_5_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4322 = io_w_req ? _GEN_3746 : CacheMem_7_5_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4323 = io_w_req ? _GEN_3747 : CacheMem_7_6_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4324 = io_w_req ? _GEN_3748 : CacheMem_7_6_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4325 = io_w_req ? _GEN_3749 : CacheMem_7_6_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4326 = io_w_req ? _GEN_3750 : CacheMem_7_6_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4327 = io_w_req ? _GEN_3751 : CacheMem_7_6_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4328 = io_w_req ? _GEN_3752 : CacheMem_7_6_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4329 = io_w_req ? _GEN_3753 : CacheMem_7_6_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4330 = io_w_req ? _GEN_3754 : CacheMem_7_6_7; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4331 = io_w_req ? _GEN_3755 : CacheMem_7_7_0; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4332 = io_w_req ? _GEN_3756 : CacheMem_7_7_1; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4333 = io_w_req ? _GEN_3757 : CacheMem_7_7_2; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4334 = io_w_req ? _GEN_3758 : CacheMem_7_7_3; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4335 = io_w_req ? _GEN_3759 : CacheMem_7_7_4; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4336 = io_w_req ? _GEN_3760 : CacheMem_7_7_5; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4337 = io_w_req ? _GEN_3761 : CacheMem_7_7_6; // @[Cache.scala 132:40 53:25]
  wire [31:0] _GEN_4338 = io_w_req ? _GEN_3762 : CacheMem_7_7_7; // @[Cache.scala 132:40 53:25]
  wire  _GEN_4339 = io_w_req ? _GEN_3763 : dirty_0_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4340 = io_w_req ? _GEN_3764 : dirty_0_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4341 = io_w_req ? _GEN_3765 : dirty_0_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4342 = io_w_req ? _GEN_3766 : dirty_0_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4343 = io_w_req ? _GEN_3767 : dirty_0_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4344 = io_w_req ? _GEN_3768 : dirty_0_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4345 = io_w_req ? _GEN_3769 : dirty_0_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4346 = io_w_req ? _GEN_3770 : dirty_0_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4347 = io_w_req ? _GEN_3771 : dirty_1_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4348 = io_w_req ? _GEN_3772 : dirty_1_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4349 = io_w_req ? _GEN_3773 : dirty_1_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4350 = io_w_req ? _GEN_3774 : dirty_1_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4351 = io_w_req ? _GEN_3775 : dirty_1_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4352 = io_w_req ? _GEN_3776 : dirty_1_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4353 = io_w_req ? _GEN_3777 : dirty_1_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4354 = io_w_req ? _GEN_3778 : dirty_1_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4355 = io_w_req ? _GEN_3779 : dirty_2_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4356 = io_w_req ? _GEN_3780 : dirty_2_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4357 = io_w_req ? _GEN_3781 : dirty_2_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4358 = io_w_req ? _GEN_3782 : dirty_2_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4359 = io_w_req ? _GEN_3783 : dirty_2_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4360 = io_w_req ? _GEN_3784 : dirty_2_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4361 = io_w_req ? _GEN_3785 : dirty_2_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4362 = io_w_req ? _GEN_3786 : dirty_2_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4363 = io_w_req ? _GEN_3787 : dirty_3_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4364 = io_w_req ? _GEN_3788 : dirty_3_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4365 = io_w_req ? _GEN_3789 : dirty_3_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4366 = io_w_req ? _GEN_3790 : dirty_3_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4367 = io_w_req ? _GEN_3791 : dirty_3_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4368 = io_w_req ? _GEN_3792 : dirty_3_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4369 = io_w_req ? _GEN_3793 : dirty_3_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4370 = io_w_req ? _GEN_3794 : dirty_3_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4371 = io_w_req ? _GEN_3795 : dirty_4_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4372 = io_w_req ? _GEN_3796 : dirty_4_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4373 = io_w_req ? _GEN_3797 : dirty_4_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4374 = io_w_req ? _GEN_3798 : dirty_4_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4375 = io_w_req ? _GEN_3799 : dirty_4_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4376 = io_w_req ? _GEN_3800 : dirty_4_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4377 = io_w_req ? _GEN_3801 : dirty_4_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4378 = io_w_req ? _GEN_3802 : dirty_4_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4379 = io_w_req ? _GEN_3803 : dirty_5_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4380 = io_w_req ? _GEN_3804 : dirty_5_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4381 = io_w_req ? _GEN_3805 : dirty_5_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4382 = io_w_req ? _GEN_3806 : dirty_5_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4383 = io_w_req ? _GEN_3807 : dirty_5_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4384 = io_w_req ? _GEN_3808 : dirty_5_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4385 = io_w_req ? _GEN_3809 : dirty_5_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4386 = io_w_req ? _GEN_3810 : dirty_5_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4387 = io_w_req ? _GEN_3811 : dirty_6_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4388 = io_w_req ? _GEN_3812 : dirty_6_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4389 = io_w_req ? _GEN_3813 : dirty_6_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4390 = io_w_req ? _GEN_3814 : dirty_6_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4391 = io_w_req ? _GEN_3815 : dirty_6_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4392 = io_w_req ? _GEN_3816 : dirty_6_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4393 = io_w_req ? _GEN_3817 : dirty_6_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4394 = io_w_req ? _GEN_3818 : dirty_6_7; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4395 = io_w_req ? _GEN_3819 : dirty_7_0; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4396 = io_w_req ? _GEN_3820 : dirty_7_1; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4397 = io_w_req ? _GEN_3821 : dirty_7_2; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4398 = io_w_req ? _GEN_3822 : dirty_7_3; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4399 = io_w_req ? _GEN_3823 : dirty_7_4; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4400 = io_w_req ? _GEN_3824 : dirty_7_5; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4401 = io_w_req ? _GEN_3825 : dirty_7_6; // @[Cache.scala 132:40 58:22]
  wire  _GEN_4402 = io_w_req ? _GEN_3826 : dirty_7_7; // @[Cache.scala 132:40 58:22]
  wire [1:0] _GEN_4403 = io_w_req ? cacheState : 2'h0; // @[Cache.scala 132:40 146:22 96:27]
  wire [31:0] _GEN_4404 = io_r_req ? _GEN_690 : 32'h0; // @[Cache.scala 129:34 131:15]
  wire [2:0] wayout_choice = _GEN_170[2:0];
  wire  _GEN_18216 = 3'h1 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4983 = _GEN_9835 & 3'h1 == wayout_choice ? valid_0_1 : valid_0_0; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18218 = 3'h2 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4984 = _GEN_9835 & 3'h2 == wayout_choice ? valid_0_2 : _GEN_4983; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18220 = 3'h3 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4985 = _GEN_9835 & 3'h3 == wayout_choice ? valid_0_3 : _GEN_4984; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18222 = 3'h4 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4986 = _GEN_9835 & 3'h4 == wayout_choice ? valid_0_4 : _GEN_4985; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18224 = 3'h5 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4987 = _GEN_9835 & 3'h5 == wayout_choice ? valid_0_5 : _GEN_4986; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18226 = 3'h6 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4988 = _GEN_9835 & 3'h6 == wayout_choice ? valid_0_6 : _GEN_4987; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18228 = 3'h7 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4989 = _GEN_9835 & 3'h7 == wayout_choice ? valid_0_7 : _GEN_4988; // @[Cache.scala 150:{47,47}]
  wire  _GEN_18230 = 3'h0 == wayout_choice; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4990 = _GEN_10087 & 3'h0 == wayout_choice ? valid_1_0 : _GEN_4989; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4991 = _GEN_10087 & 3'h1 == wayout_choice ? valid_1_1 : _GEN_4990; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4992 = _GEN_10087 & 3'h2 == wayout_choice ? valid_1_2 : _GEN_4991; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4993 = _GEN_10087 & 3'h3 == wayout_choice ? valid_1_3 : _GEN_4992; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4994 = _GEN_10087 & 3'h4 == wayout_choice ? valid_1_4 : _GEN_4993; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4995 = _GEN_10087 & 3'h5 == wayout_choice ? valid_1_5 : _GEN_4994; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4996 = _GEN_10087 & 3'h6 == wayout_choice ? valid_1_6 : _GEN_4995; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4997 = _GEN_10087 & 3'h7 == wayout_choice ? valid_1_7 : _GEN_4996; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4998 = _GEN_10343 & 3'h0 == wayout_choice ? valid_2_0 : _GEN_4997; // @[Cache.scala 150:{47,47}]
  wire  _GEN_4999 = _GEN_10343 & 3'h1 == wayout_choice ? valid_2_1 : _GEN_4998; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5000 = _GEN_10343 & 3'h2 == wayout_choice ? valid_2_2 : _GEN_4999; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5001 = _GEN_10343 & 3'h3 == wayout_choice ? valid_2_3 : _GEN_5000; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5002 = _GEN_10343 & 3'h4 == wayout_choice ? valid_2_4 : _GEN_5001; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5003 = _GEN_10343 & 3'h5 == wayout_choice ? valid_2_5 : _GEN_5002; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5004 = _GEN_10343 & 3'h6 == wayout_choice ? valid_2_6 : _GEN_5003; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5005 = _GEN_10343 & 3'h7 == wayout_choice ? valid_2_7 : _GEN_5004; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5006 = _GEN_10599 & 3'h0 == wayout_choice ? valid_3_0 : _GEN_5005; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5007 = _GEN_10599 & 3'h1 == wayout_choice ? valid_3_1 : _GEN_5006; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5008 = _GEN_10599 & 3'h2 == wayout_choice ? valid_3_2 : _GEN_5007; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5009 = _GEN_10599 & 3'h3 == wayout_choice ? valid_3_3 : _GEN_5008; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5010 = _GEN_10599 & 3'h4 == wayout_choice ? valid_3_4 : _GEN_5009; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5011 = _GEN_10599 & 3'h5 == wayout_choice ? valid_3_5 : _GEN_5010; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5012 = _GEN_10599 & 3'h6 == wayout_choice ? valid_3_6 : _GEN_5011; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5013 = _GEN_10599 & 3'h7 == wayout_choice ? valid_3_7 : _GEN_5012; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5014 = _GEN_10855 & 3'h0 == wayout_choice ? valid_4_0 : _GEN_5013; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5015 = _GEN_10855 & 3'h1 == wayout_choice ? valid_4_1 : _GEN_5014; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5016 = _GEN_10855 & 3'h2 == wayout_choice ? valid_4_2 : _GEN_5015; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5017 = _GEN_10855 & 3'h3 == wayout_choice ? valid_4_3 : _GEN_5016; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5018 = _GEN_10855 & 3'h4 == wayout_choice ? valid_4_4 : _GEN_5017; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5019 = _GEN_10855 & 3'h5 == wayout_choice ? valid_4_5 : _GEN_5018; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5020 = _GEN_10855 & 3'h6 == wayout_choice ? valid_4_6 : _GEN_5019; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5021 = _GEN_10855 & 3'h7 == wayout_choice ? valid_4_7 : _GEN_5020; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5022 = _GEN_11111 & 3'h0 == wayout_choice ? valid_5_0 : _GEN_5021; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5023 = _GEN_11111 & 3'h1 == wayout_choice ? valid_5_1 : _GEN_5022; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5024 = _GEN_11111 & 3'h2 == wayout_choice ? valid_5_2 : _GEN_5023; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5025 = _GEN_11111 & 3'h3 == wayout_choice ? valid_5_3 : _GEN_5024; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5026 = _GEN_11111 & 3'h4 == wayout_choice ? valid_5_4 : _GEN_5025; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5027 = _GEN_11111 & 3'h5 == wayout_choice ? valid_5_5 : _GEN_5026; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5028 = _GEN_11111 & 3'h6 == wayout_choice ? valid_5_6 : _GEN_5027; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5029 = _GEN_11111 & 3'h7 == wayout_choice ? valid_5_7 : _GEN_5028; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5030 = _GEN_11367 & 3'h0 == wayout_choice ? valid_6_0 : _GEN_5029; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5031 = _GEN_11367 & 3'h1 == wayout_choice ? valid_6_1 : _GEN_5030; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5032 = _GEN_11367 & 3'h2 == wayout_choice ? valid_6_2 : _GEN_5031; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5033 = _GEN_11367 & 3'h3 == wayout_choice ? valid_6_3 : _GEN_5032; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5034 = _GEN_11367 & 3'h4 == wayout_choice ? valid_6_4 : _GEN_5033; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5035 = _GEN_11367 & 3'h5 == wayout_choice ? valid_6_5 : _GEN_5034; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5036 = _GEN_11367 & 3'h6 == wayout_choice ? valid_6_6 : _GEN_5035; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5037 = _GEN_11367 & 3'h7 == wayout_choice ? valid_6_7 : _GEN_5036; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5038 = _GEN_11623 & 3'h0 == wayout_choice ? valid_7_0 : _GEN_5037; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5039 = _GEN_11623 & 3'h1 == wayout_choice ? valid_7_1 : _GEN_5038; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5040 = _GEN_11623 & 3'h2 == wayout_choice ? valid_7_2 : _GEN_5039; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5041 = _GEN_11623 & 3'h3 == wayout_choice ? valid_7_3 : _GEN_5040; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5042 = _GEN_11623 & 3'h4 == wayout_choice ? valid_7_4 : _GEN_5041; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5043 = _GEN_11623 & 3'h5 == wayout_choice ? valid_7_5 : _GEN_5042; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5044 = _GEN_11623 & 3'h6 == wayout_choice ? valid_7_6 : _GEN_5043; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5045 = _GEN_11623 & 3'h7 == wayout_choice ? valid_7_7 : _GEN_5044; // @[Cache.scala 150:{47,47}]
  wire  _GEN_5047 = _GEN_9835 & 3'h1 == wayout_choice ? dirty_0_1 : dirty_0_0; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5048 = _GEN_9835 & 3'h2 == wayout_choice ? dirty_0_2 : _GEN_5047; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5049 = _GEN_9835 & 3'h3 == wayout_choice ? dirty_0_3 : _GEN_5048; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5050 = _GEN_9835 & 3'h4 == wayout_choice ? dirty_0_4 : _GEN_5049; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5051 = _GEN_9835 & 3'h5 == wayout_choice ? dirty_0_5 : _GEN_5050; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5052 = _GEN_9835 & 3'h6 == wayout_choice ? dirty_0_6 : _GEN_5051; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5053 = _GEN_9835 & 3'h7 == wayout_choice ? dirty_0_7 : _GEN_5052; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5054 = _GEN_10087 & 3'h0 == wayout_choice ? dirty_1_0 : _GEN_5053; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5055 = _GEN_10087 & 3'h1 == wayout_choice ? dirty_1_1 : _GEN_5054; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5056 = _GEN_10087 & 3'h2 == wayout_choice ? dirty_1_2 : _GEN_5055; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5057 = _GEN_10087 & 3'h3 == wayout_choice ? dirty_1_3 : _GEN_5056; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5058 = _GEN_10087 & 3'h4 == wayout_choice ? dirty_1_4 : _GEN_5057; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5059 = _GEN_10087 & 3'h5 == wayout_choice ? dirty_1_5 : _GEN_5058; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5060 = _GEN_10087 & 3'h6 == wayout_choice ? dirty_1_6 : _GEN_5059; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5061 = _GEN_10087 & 3'h7 == wayout_choice ? dirty_1_7 : _GEN_5060; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5062 = _GEN_10343 & 3'h0 == wayout_choice ? dirty_2_0 : _GEN_5061; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5063 = _GEN_10343 & 3'h1 == wayout_choice ? dirty_2_1 : _GEN_5062; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5064 = _GEN_10343 & 3'h2 == wayout_choice ? dirty_2_2 : _GEN_5063; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5065 = _GEN_10343 & 3'h3 == wayout_choice ? dirty_2_3 : _GEN_5064; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5066 = _GEN_10343 & 3'h4 == wayout_choice ? dirty_2_4 : _GEN_5065; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5067 = _GEN_10343 & 3'h5 == wayout_choice ? dirty_2_5 : _GEN_5066; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5068 = _GEN_10343 & 3'h6 == wayout_choice ? dirty_2_6 : _GEN_5067; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5069 = _GEN_10343 & 3'h7 == wayout_choice ? dirty_2_7 : _GEN_5068; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5070 = _GEN_10599 & 3'h0 == wayout_choice ? dirty_3_0 : _GEN_5069; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5071 = _GEN_10599 & 3'h1 == wayout_choice ? dirty_3_1 : _GEN_5070; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5072 = _GEN_10599 & 3'h2 == wayout_choice ? dirty_3_2 : _GEN_5071; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5073 = _GEN_10599 & 3'h3 == wayout_choice ? dirty_3_3 : _GEN_5072; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5074 = _GEN_10599 & 3'h4 == wayout_choice ? dirty_3_4 : _GEN_5073; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5075 = _GEN_10599 & 3'h5 == wayout_choice ? dirty_3_5 : _GEN_5074; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5076 = _GEN_10599 & 3'h6 == wayout_choice ? dirty_3_6 : _GEN_5075; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5077 = _GEN_10599 & 3'h7 == wayout_choice ? dirty_3_7 : _GEN_5076; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5078 = _GEN_10855 & 3'h0 == wayout_choice ? dirty_4_0 : _GEN_5077; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5079 = _GEN_10855 & 3'h1 == wayout_choice ? dirty_4_1 : _GEN_5078; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5080 = _GEN_10855 & 3'h2 == wayout_choice ? dirty_4_2 : _GEN_5079; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5081 = _GEN_10855 & 3'h3 == wayout_choice ? dirty_4_3 : _GEN_5080; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5082 = _GEN_10855 & 3'h4 == wayout_choice ? dirty_4_4 : _GEN_5081; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5083 = _GEN_10855 & 3'h5 == wayout_choice ? dirty_4_5 : _GEN_5082; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5084 = _GEN_10855 & 3'h6 == wayout_choice ? dirty_4_6 : _GEN_5083; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5085 = _GEN_10855 & 3'h7 == wayout_choice ? dirty_4_7 : _GEN_5084; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5086 = _GEN_11111 & 3'h0 == wayout_choice ? dirty_5_0 : _GEN_5085; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5087 = _GEN_11111 & 3'h1 == wayout_choice ? dirty_5_1 : _GEN_5086; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5088 = _GEN_11111 & 3'h2 == wayout_choice ? dirty_5_2 : _GEN_5087; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5089 = _GEN_11111 & 3'h3 == wayout_choice ? dirty_5_3 : _GEN_5088; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5090 = _GEN_11111 & 3'h4 == wayout_choice ? dirty_5_4 : _GEN_5089; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5091 = _GEN_11111 & 3'h5 == wayout_choice ? dirty_5_5 : _GEN_5090; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5092 = _GEN_11111 & 3'h6 == wayout_choice ? dirty_5_6 : _GEN_5091; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5093 = _GEN_11111 & 3'h7 == wayout_choice ? dirty_5_7 : _GEN_5092; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5094 = _GEN_11367 & 3'h0 == wayout_choice ? dirty_6_0 : _GEN_5093; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5095 = _GEN_11367 & 3'h1 == wayout_choice ? dirty_6_1 : _GEN_5094; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5096 = _GEN_11367 & 3'h2 == wayout_choice ? dirty_6_2 : _GEN_5095; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5097 = _GEN_11367 & 3'h3 == wayout_choice ? dirty_6_3 : _GEN_5096; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5098 = _GEN_11367 & 3'h4 == wayout_choice ? dirty_6_4 : _GEN_5097; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5099 = _GEN_11367 & 3'h5 == wayout_choice ? dirty_6_5 : _GEN_5098; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5100 = _GEN_11367 & 3'h6 == wayout_choice ? dirty_6_6 : _GEN_5099; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5101 = _GEN_11367 & 3'h7 == wayout_choice ? dirty_6_7 : _GEN_5100; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5102 = _GEN_11623 & 3'h0 == wayout_choice ? dirty_7_0 : _GEN_5101; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5103 = _GEN_11623 & 3'h1 == wayout_choice ? dirty_7_1 : _GEN_5102; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5104 = _GEN_11623 & 3'h2 == wayout_choice ? dirty_7_2 : _GEN_5103; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5105 = _GEN_11623 & 3'h3 == wayout_choice ? dirty_7_3 : _GEN_5104; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5106 = _GEN_11623 & 3'h4 == wayout_choice ? dirty_7_4 : _GEN_5105; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5107 = _GEN_11623 & 3'h5 == wayout_choice ? dirty_7_5 : _GEN_5106; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5108 = _GEN_11623 & 3'h6 == wayout_choice ? dirty_7_6 : _GEN_5107; // @[Cache.scala 150:{92,92}]
  wire  _GEN_5109 = _GEN_11623 & 3'h7 == wayout_choice ? dirty_7_7 : _GEN_5108; // @[Cache.scala 150:{92,92}]
  wire [5:0] _GEN_5111 = _GEN_9835 & _GEN_18216 ? cache_tags_0_1 : cache_tags_0_0; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5112 = _GEN_9835 & _GEN_18218 ? cache_tags_0_2 : _GEN_5111; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5113 = _GEN_9835 & _GEN_18220 ? cache_tags_0_3 : _GEN_5112; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5114 = _GEN_9835 & _GEN_18222 ? cache_tags_0_4 : _GEN_5113; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5115 = _GEN_9835 & _GEN_18224 ? cache_tags_0_5 : _GEN_5114; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5116 = _GEN_9835 & _GEN_18226 ? cache_tags_0_6 : _GEN_5115; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5117 = _GEN_9835 & _GEN_18228 ? cache_tags_0_7 : _GEN_5116; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5118 = _GEN_10087 & _GEN_18230 ? cache_tags_1_0 : _GEN_5117; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5119 = _GEN_10087 & _GEN_18216 ? cache_tags_1_1 : _GEN_5118; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5120 = _GEN_10087 & _GEN_18218 ? cache_tags_1_2 : _GEN_5119; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5121 = _GEN_10087 & _GEN_18220 ? cache_tags_1_3 : _GEN_5120; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5122 = _GEN_10087 & _GEN_18222 ? cache_tags_1_4 : _GEN_5121; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5123 = _GEN_10087 & _GEN_18224 ? cache_tags_1_5 : _GEN_5122; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5124 = _GEN_10087 & _GEN_18226 ? cache_tags_1_6 : _GEN_5123; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5125 = _GEN_10087 & _GEN_18228 ? cache_tags_1_7 : _GEN_5124; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5126 = _GEN_10343 & _GEN_18230 ? cache_tags_2_0 : _GEN_5125; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5127 = _GEN_10343 & _GEN_18216 ? cache_tags_2_1 : _GEN_5126; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5128 = _GEN_10343 & _GEN_18218 ? cache_tags_2_2 : _GEN_5127; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5129 = _GEN_10343 & _GEN_18220 ? cache_tags_2_3 : _GEN_5128; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5130 = _GEN_10343 & _GEN_18222 ? cache_tags_2_4 : _GEN_5129; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5131 = _GEN_10343 & _GEN_18224 ? cache_tags_2_5 : _GEN_5130; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5132 = _GEN_10343 & _GEN_18226 ? cache_tags_2_6 : _GEN_5131; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5133 = _GEN_10343 & _GEN_18228 ? cache_tags_2_7 : _GEN_5132; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5134 = _GEN_10599 & _GEN_18230 ? cache_tags_3_0 : _GEN_5133; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5135 = _GEN_10599 & _GEN_18216 ? cache_tags_3_1 : _GEN_5134; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5136 = _GEN_10599 & _GEN_18218 ? cache_tags_3_2 : _GEN_5135; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5137 = _GEN_10599 & _GEN_18220 ? cache_tags_3_3 : _GEN_5136; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5138 = _GEN_10599 & _GEN_18222 ? cache_tags_3_4 : _GEN_5137; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5139 = _GEN_10599 & _GEN_18224 ? cache_tags_3_5 : _GEN_5138; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5140 = _GEN_10599 & _GEN_18226 ? cache_tags_3_6 : _GEN_5139; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5141 = _GEN_10599 & _GEN_18228 ? cache_tags_3_7 : _GEN_5140; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5142 = _GEN_10855 & _GEN_18230 ? cache_tags_4_0 : _GEN_5141; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5143 = _GEN_10855 & _GEN_18216 ? cache_tags_4_1 : _GEN_5142; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5144 = _GEN_10855 & _GEN_18218 ? cache_tags_4_2 : _GEN_5143; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5145 = _GEN_10855 & _GEN_18220 ? cache_tags_4_3 : _GEN_5144; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5146 = _GEN_10855 & _GEN_18222 ? cache_tags_4_4 : _GEN_5145; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5147 = _GEN_10855 & _GEN_18224 ? cache_tags_4_5 : _GEN_5146; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5148 = _GEN_10855 & _GEN_18226 ? cache_tags_4_6 : _GEN_5147; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5149 = _GEN_10855 & _GEN_18228 ? cache_tags_4_7 : _GEN_5148; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5150 = _GEN_11111 & _GEN_18230 ? cache_tags_5_0 : _GEN_5149; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5151 = _GEN_11111 & _GEN_18216 ? cache_tags_5_1 : _GEN_5150; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5152 = _GEN_11111 & _GEN_18218 ? cache_tags_5_2 : _GEN_5151; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5153 = _GEN_11111 & _GEN_18220 ? cache_tags_5_3 : _GEN_5152; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5154 = _GEN_11111 & _GEN_18222 ? cache_tags_5_4 : _GEN_5153; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5155 = _GEN_11111 & _GEN_18224 ? cache_tags_5_5 : _GEN_5154; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5156 = _GEN_11111 & _GEN_18226 ? cache_tags_5_6 : _GEN_5155; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5157 = _GEN_11111 & _GEN_18228 ? cache_tags_5_7 : _GEN_5156; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5158 = _GEN_11367 & _GEN_18230 ? cache_tags_6_0 : _GEN_5157; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5159 = _GEN_11367 & _GEN_18216 ? cache_tags_6_1 : _GEN_5158; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5160 = _GEN_11367 & _GEN_18218 ? cache_tags_6_2 : _GEN_5159; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5161 = _GEN_11367 & _GEN_18220 ? cache_tags_6_3 : _GEN_5160; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5162 = _GEN_11367 & _GEN_18222 ? cache_tags_6_4 : _GEN_5161; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5163 = _GEN_11367 & _GEN_18224 ? cache_tags_6_5 : _GEN_5162; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5164 = _GEN_11367 & _GEN_18226 ? cache_tags_6_6 : _GEN_5163; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5165 = _GEN_11367 & _GEN_18228 ? cache_tags_6_7 : _GEN_5164; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5166 = _GEN_11623 & _GEN_18230 ? cache_tags_7_0 : _GEN_5165; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5167 = _GEN_11623 & _GEN_18216 ? cache_tags_7_1 : _GEN_5166; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5168 = _GEN_11623 & _GEN_18218 ? cache_tags_7_2 : _GEN_5167; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5169 = _GEN_11623 & _GEN_18220 ? cache_tags_7_3 : _GEN_5168; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5170 = _GEN_11623 & _GEN_18222 ? cache_tags_7_4 : _GEN_5169; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5171 = _GEN_11623 & _GEN_18224 ? cache_tags_7_5 : _GEN_5170; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5172 = _GEN_11623 & _GEN_18226 ? cache_tags_7_6 : _GEN_5171; // @[Cat.scala 31:{58,58}]
  wire [5:0] _GEN_5173 = _GEN_11623 & _GEN_18228 ? cache_tags_7_7 : _GEN_5172; // @[Cat.scala 31:{58,58}]
  wire [8:0] _mem_wr_addr_T = {_GEN_5173,set_addr}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_5175 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_0 : CacheMem_0_0_0; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5176 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_0 : _GEN_5175; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5177 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_0 : _GEN_5176; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5178 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_0 : _GEN_5177; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5179 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_0 : _GEN_5178; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5180 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_0 : _GEN_5179; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5181 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_0 : _GEN_5180; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5182 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_0 : _GEN_5181; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5183 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_0 : _GEN_5182; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5184 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_0 : _GEN_5183; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5185 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_0 : _GEN_5184; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5186 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_0 : _GEN_5185; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5187 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_0 : _GEN_5186; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5188 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_0 : _GEN_5187; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5189 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_0 : _GEN_5188; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5190 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_0 : _GEN_5189; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5191 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_0 : _GEN_5190; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5192 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_0 : _GEN_5191; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5193 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_0 : _GEN_5192; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5194 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_0 : _GEN_5193; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5195 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_0 : _GEN_5194; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5196 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_0 : _GEN_5195; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5197 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_0 : _GEN_5196; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5198 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_0 : _GEN_5197; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5199 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_0 : _GEN_5198; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5200 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_0 : _GEN_5199; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5201 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_0 : _GEN_5200; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5202 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_0 : _GEN_5201; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5203 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_0 : _GEN_5202; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5204 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_0 : _GEN_5203; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5205 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_0 : _GEN_5204; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5206 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_0 : _GEN_5205; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5207 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_0 : _GEN_5206; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5208 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_0 : _GEN_5207; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5209 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_0 : _GEN_5208; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5210 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_0 : _GEN_5209; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5211 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_0 : _GEN_5210; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5212 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_0 : _GEN_5211; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5213 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_0 : _GEN_5212; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5214 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_0 : _GEN_5213; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5215 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_0 : _GEN_5214; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5216 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_0 : _GEN_5215; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5217 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_0 : _GEN_5216; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5218 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_0 : _GEN_5217; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5219 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_0 : _GEN_5218; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5220 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_0 : _GEN_5219; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5221 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_0 : _GEN_5220; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5222 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_0 : _GEN_5221; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5223 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_0 : _GEN_5222; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5224 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_0 : _GEN_5223; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5225 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_0 : _GEN_5224; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5226 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_0 : _GEN_5225; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5227 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_0 : _GEN_5226; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5228 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_0 : _GEN_5227; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5229 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_0 : _GEN_5228; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5230 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_0 : _GEN_5229; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5231 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_0 : _GEN_5230; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5232 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_0 : _GEN_5231; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5233 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_0 : _GEN_5232; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5234 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_0 : _GEN_5233; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5235 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_0 : _GEN_5234; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5236 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_0 : _GEN_5235; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5237 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_0 : _GEN_5236; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5239 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_1 : CacheMem_0_0_1; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5240 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_1 : _GEN_5239; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5241 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_1 : _GEN_5240; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5242 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_1 : _GEN_5241; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5243 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_1 : _GEN_5242; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5244 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_1 : _GEN_5243; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5245 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_1 : _GEN_5244; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5246 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_1 : _GEN_5245; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5247 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_1 : _GEN_5246; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5248 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_1 : _GEN_5247; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5249 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_1 : _GEN_5248; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5250 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_1 : _GEN_5249; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5251 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_1 : _GEN_5250; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5252 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_1 : _GEN_5251; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5253 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_1 : _GEN_5252; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5254 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_1 : _GEN_5253; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5255 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_1 : _GEN_5254; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5256 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_1 : _GEN_5255; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5257 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_1 : _GEN_5256; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5258 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_1 : _GEN_5257; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5259 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_1 : _GEN_5258; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5260 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_1 : _GEN_5259; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5261 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_1 : _GEN_5260; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5262 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_1 : _GEN_5261; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5263 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_1 : _GEN_5262; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5264 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_1 : _GEN_5263; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5265 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_1 : _GEN_5264; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5266 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_1 : _GEN_5265; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5267 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_1 : _GEN_5266; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5268 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_1 : _GEN_5267; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5269 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_1 : _GEN_5268; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5270 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_1 : _GEN_5269; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5271 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_1 : _GEN_5270; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5272 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_1 : _GEN_5271; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5273 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_1 : _GEN_5272; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5274 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_1 : _GEN_5273; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5275 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_1 : _GEN_5274; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5276 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_1 : _GEN_5275; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5277 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_1 : _GEN_5276; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5278 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_1 : _GEN_5277; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5279 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_1 : _GEN_5278; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5280 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_1 : _GEN_5279; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5281 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_1 : _GEN_5280; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5282 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_1 : _GEN_5281; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5283 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_1 : _GEN_5282; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5284 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_1 : _GEN_5283; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5285 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_1 : _GEN_5284; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5286 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_1 : _GEN_5285; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5287 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_1 : _GEN_5286; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5288 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_1 : _GEN_5287; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5289 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_1 : _GEN_5288; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5290 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_1 : _GEN_5289; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5291 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_1 : _GEN_5290; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5292 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_1 : _GEN_5291; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5293 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_1 : _GEN_5292; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5294 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_1 : _GEN_5293; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5295 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_1 : _GEN_5294; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5296 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_1 : _GEN_5295; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5297 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_1 : _GEN_5296; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5298 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_1 : _GEN_5297; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5299 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_1 : _GEN_5298; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5300 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_1 : _GEN_5299; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5301 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_1 : _GEN_5300; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5303 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_2 : CacheMem_0_0_2; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5304 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_2 : _GEN_5303; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5305 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_2 : _GEN_5304; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5306 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_2 : _GEN_5305; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5307 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_2 : _GEN_5306; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5308 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_2 : _GEN_5307; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5309 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_2 : _GEN_5308; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5310 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_2 : _GEN_5309; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5311 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_2 : _GEN_5310; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5312 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_2 : _GEN_5311; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5313 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_2 : _GEN_5312; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5314 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_2 : _GEN_5313; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5315 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_2 : _GEN_5314; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5316 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_2 : _GEN_5315; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5317 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_2 : _GEN_5316; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5318 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_2 : _GEN_5317; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5319 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_2 : _GEN_5318; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5320 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_2 : _GEN_5319; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5321 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_2 : _GEN_5320; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5322 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_2 : _GEN_5321; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5323 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_2 : _GEN_5322; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5324 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_2 : _GEN_5323; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5325 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_2 : _GEN_5324; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5326 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_2 : _GEN_5325; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5327 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_2 : _GEN_5326; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5328 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_2 : _GEN_5327; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5329 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_2 : _GEN_5328; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5330 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_2 : _GEN_5329; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5331 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_2 : _GEN_5330; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5332 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_2 : _GEN_5331; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5333 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_2 : _GEN_5332; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5334 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_2 : _GEN_5333; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5335 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_2 : _GEN_5334; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5336 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_2 : _GEN_5335; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5337 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_2 : _GEN_5336; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5338 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_2 : _GEN_5337; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5339 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_2 : _GEN_5338; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5340 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_2 : _GEN_5339; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5341 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_2 : _GEN_5340; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5342 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_2 : _GEN_5341; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5343 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_2 : _GEN_5342; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5344 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_2 : _GEN_5343; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5345 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_2 : _GEN_5344; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5346 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_2 : _GEN_5345; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5347 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_2 : _GEN_5346; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5348 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_2 : _GEN_5347; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5349 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_2 : _GEN_5348; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5350 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_2 : _GEN_5349; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5351 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_2 : _GEN_5350; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5352 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_2 : _GEN_5351; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5353 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_2 : _GEN_5352; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5354 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_2 : _GEN_5353; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5355 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_2 : _GEN_5354; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5356 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_2 : _GEN_5355; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5357 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_2 : _GEN_5356; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5358 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_2 : _GEN_5357; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5359 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_2 : _GEN_5358; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5360 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_2 : _GEN_5359; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5361 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_2 : _GEN_5360; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5362 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_2 : _GEN_5361; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5363 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_2 : _GEN_5362; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5364 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_2 : _GEN_5363; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5365 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_2 : _GEN_5364; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5367 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_3 : CacheMem_0_0_3; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5368 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_3 : _GEN_5367; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5369 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_3 : _GEN_5368; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5370 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_3 : _GEN_5369; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5371 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_3 : _GEN_5370; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5372 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_3 : _GEN_5371; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5373 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_3 : _GEN_5372; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5374 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_3 : _GEN_5373; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5375 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_3 : _GEN_5374; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5376 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_3 : _GEN_5375; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5377 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_3 : _GEN_5376; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5378 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_3 : _GEN_5377; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5379 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_3 : _GEN_5378; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5380 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_3 : _GEN_5379; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5381 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_3 : _GEN_5380; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5382 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_3 : _GEN_5381; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5383 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_3 : _GEN_5382; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5384 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_3 : _GEN_5383; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5385 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_3 : _GEN_5384; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5386 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_3 : _GEN_5385; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5387 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_3 : _GEN_5386; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5388 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_3 : _GEN_5387; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5389 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_3 : _GEN_5388; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5390 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_3 : _GEN_5389; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5391 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_3 : _GEN_5390; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5392 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_3 : _GEN_5391; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5393 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_3 : _GEN_5392; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5394 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_3 : _GEN_5393; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5395 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_3 : _GEN_5394; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5396 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_3 : _GEN_5395; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5397 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_3 : _GEN_5396; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5398 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_3 : _GEN_5397; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5399 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_3 : _GEN_5398; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5400 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_3 : _GEN_5399; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5401 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_3 : _GEN_5400; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5402 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_3 : _GEN_5401; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5403 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_3 : _GEN_5402; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5404 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_3 : _GEN_5403; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5405 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_3 : _GEN_5404; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5406 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_3 : _GEN_5405; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5407 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_3 : _GEN_5406; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5408 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_3 : _GEN_5407; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5409 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_3 : _GEN_5408; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5410 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_3 : _GEN_5409; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5411 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_3 : _GEN_5410; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5412 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_3 : _GEN_5411; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5413 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_3 : _GEN_5412; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5414 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_3 : _GEN_5413; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5415 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_3 : _GEN_5414; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5416 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_3 : _GEN_5415; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5417 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_3 : _GEN_5416; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5418 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_3 : _GEN_5417; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5419 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_3 : _GEN_5418; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5420 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_3 : _GEN_5419; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5421 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_3 : _GEN_5420; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5422 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_3 : _GEN_5421; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5423 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_3 : _GEN_5422; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5424 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_3 : _GEN_5423; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5425 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_3 : _GEN_5424; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5426 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_3 : _GEN_5425; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5427 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_3 : _GEN_5426; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5428 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_3 : _GEN_5427; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5429 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_3 : _GEN_5428; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5431 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_4 : CacheMem_0_0_4; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5432 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_4 : _GEN_5431; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5433 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_4 : _GEN_5432; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5434 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_4 : _GEN_5433; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5435 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_4 : _GEN_5434; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5436 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_4 : _GEN_5435; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5437 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_4 : _GEN_5436; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5438 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_4 : _GEN_5437; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5439 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_4 : _GEN_5438; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5440 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_4 : _GEN_5439; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5441 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_4 : _GEN_5440; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5442 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_4 : _GEN_5441; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5443 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_4 : _GEN_5442; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5444 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_4 : _GEN_5443; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5445 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_4 : _GEN_5444; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5446 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_4 : _GEN_5445; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5447 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_4 : _GEN_5446; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5448 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_4 : _GEN_5447; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5449 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_4 : _GEN_5448; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5450 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_4 : _GEN_5449; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5451 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_4 : _GEN_5450; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5452 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_4 : _GEN_5451; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5453 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_4 : _GEN_5452; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5454 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_4 : _GEN_5453; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5455 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_4 : _GEN_5454; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5456 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_4 : _GEN_5455; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5457 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_4 : _GEN_5456; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5458 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_4 : _GEN_5457; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5459 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_4 : _GEN_5458; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5460 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_4 : _GEN_5459; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5461 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_4 : _GEN_5460; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5462 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_4 : _GEN_5461; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5463 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_4 : _GEN_5462; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5464 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_4 : _GEN_5463; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5465 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_4 : _GEN_5464; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5466 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_4 : _GEN_5465; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5467 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_4 : _GEN_5466; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5468 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_4 : _GEN_5467; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5469 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_4 : _GEN_5468; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5470 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_4 : _GEN_5469; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5471 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_4 : _GEN_5470; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5472 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_4 : _GEN_5471; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5473 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_4 : _GEN_5472; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5474 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_4 : _GEN_5473; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5475 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_4 : _GEN_5474; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5476 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_4 : _GEN_5475; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5477 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_4 : _GEN_5476; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5478 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_4 : _GEN_5477; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5479 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_4 : _GEN_5478; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5480 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_4 : _GEN_5479; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5481 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_4 : _GEN_5480; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5482 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_4 : _GEN_5481; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5483 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_4 : _GEN_5482; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5484 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_4 : _GEN_5483; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5485 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_4 : _GEN_5484; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5486 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_4 : _GEN_5485; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5487 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_4 : _GEN_5486; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5488 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_4 : _GEN_5487; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5489 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_4 : _GEN_5488; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5490 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_4 : _GEN_5489; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5491 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_4 : _GEN_5490; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5492 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_4 : _GEN_5491; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5493 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_4 : _GEN_5492; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5495 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_5 : CacheMem_0_0_5; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5496 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_5 : _GEN_5495; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5497 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_5 : _GEN_5496; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5498 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_5 : _GEN_5497; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5499 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_5 : _GEN_5498; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5500 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_5 : _GEN_5499; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5501 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_5 : _GEN_5500; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5502 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_5 : _GEN_5501; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5503 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_5 : _GEN_5502; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5504 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_5 : _GEN_5503; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5505 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_5 : _GEN_5504; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5506 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_5 : _GEN_5505; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5507 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_5 : _GEN_5506; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5508 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_5 : _GEN_5507; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5509 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_5 : _GEN_5508; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5510 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_5 : _GEN_5509; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5511 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_5 : _GEN_5510; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5512 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_5 : _GEN_5511; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5513 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_5 : _GEN_5512; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5514 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_5 : _GEN_5513; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5515 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_5 : _GEN_5514; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5516 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_5 : _GEN_5515; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5517 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_5 : _GEN_5516; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5518 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_5 : _GEN_5517; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5519 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_5 : _GEN_5518; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5520 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_5 : _GEN_5519; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5521 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_5 : _GEN_5520; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5522 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_5 : _GEN_5521; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5523 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_5 : _GEN_5522; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5524 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_5 : _GEN_5523; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5525 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_5 : _GEN_5524; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5526 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_5 : _GEN_5525; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5527 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_5 : _GEN_5526; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5528 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_5 : _GEN_5527; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5529 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_5 : _GEN_5528; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5530 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_5 : _GEN_5529; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5531 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_5 : _GEN_5530; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5532 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_5 : _GEN_5531; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5533 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_5 : _GEN_5532; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5534 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_5 : _GEN_5533; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5535 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_5 : _GEN_5534; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5536 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_5 : _GEN_5535; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5537 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_5 : _GEN_5536; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5538 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_5 : _GEN_5537; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5539 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_5 : _GEN_5538; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5540 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_5 : _GEN_5539; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5541 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_5 : _GEN_5540; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5542 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_5 : _GEN_5541; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5543 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_5 : _GEN_5542; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5544 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_5 : _GEN_5543; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5545 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_5 : _GEN_5544; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5546 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_5 : _GEN_5545; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5547 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_5 : _GEN_5546; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5548 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_5 : _GEN_5547; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5549 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_5 : _GEN_5548; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5550 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_5 : _GEN_5549; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5551 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_5 : _GEN_5550; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5552 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_5 : _GEN_5551; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5553 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_5 : _GEN_5552; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5554 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_5 : _GEN_5553; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5555 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_5 : _GEN_5554; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5556 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_5 : _GEN_5555; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5557 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_5 : _GEN_5556; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5559 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_6 : CacheMem_0_0_6; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5560 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_6 : _GEN_5559; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5561 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_6 : _GEN_5560; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5562 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_6 : _GEN_5561; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5563 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_6 : _GEN_5562; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5564 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_6 : _GEN_5563; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5565 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_6 : _GEN_5564; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5566 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_6 : _GEN_5565; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5567 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_6 : _GEN_5566; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5568 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_6 : _GEN_5567; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5569 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_6 : _GEN_5568; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5570 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_6 : _GEN_5569; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5571 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_6 : _GEN_5570; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5572 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_6 : _GEN_5571; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5573 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_6 : _GEN_5572; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5574 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_6 : _GEN_5573; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5575 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_6 : _GEN_5574; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5576 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_6 : _GEN_5575; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5577 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_6 : _GEN_5576; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5578 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_6 : _GEN_5577; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5579 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_6 : _GEN_5578; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5580 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_6 : _GEN_5579; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5581 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_6 : _GEN_5580; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5582 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_6 : _GEN_5581; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5583 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_6 : _GEN_5582; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5584 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_6 : _GEN_5583; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5585 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_6 : _GEN_5584; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5586 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_6 : _GEN_5585; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5587 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_6 : _GEN_5586; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5588 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_6 : _GEN_5587; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5589 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_6 : _GEN_5588; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5590 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_6 : _GEN_5589; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5591 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_6 : _GEN_5590; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5592 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_6 : _GEN_5591; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5593 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_6 : _GEN_5592; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5594 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_6 : _GEN_5593; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5595 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_6 : _GEN_5594; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5596 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_6 : _GEN_5595; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5597 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_6 : _GEN_5596; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5598 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_6 : _GEN_5597; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5599 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_6 : _GEN_5598; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5600 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_6 : _GEN_5599; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5601 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_6 : _GEN_5600; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5602 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_6 : _GEN_5601; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5603 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_6 : _GEN_5602; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5604 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_6 : _GEN_5603; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5605 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_6 : _GEN_5604; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5606 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_6 : _GEN_5605; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5607 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_6 : _GEN_5606; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5608 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_6 : _GEN_5607; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5609 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_6 : _GEN_5608; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5610 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_6 : _GEN_5609; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5611 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_6 : _GEN_5610; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5612 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_6 : _GEN_5611; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5613 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_6 : _GEN_5612; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5614 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_6 : _GEN_5613; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5615 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_6 : _GEN_5614; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5616 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_6 : _GEN_5615; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5617 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_6 : _GEN_5616; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5618 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_6 : _GEN_5617; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5619 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_6 : _GEN_5618; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5620 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_6 : _GEN_5619; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5621 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_6 : _GEN_5620; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5623 = _GEN_9835 & _GEN_18216 ? CacheMem_0_1_7 : CacheMem_0_0_7; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5624 = _GEN_9835 & _GEN_18218 ? CacheMem_0_2_7 : _GEN_5623; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5625 = _GEN_9835 & _GEN_18220 ? CacheMem_0_3_7 : _GEN_5624; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5626 = _GEN_9835 & _GEN_18222 ? CacheMem_0_4_7 : _GEN_5625; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5627 = _GEN_9835 & _GEN_18224 ? CacheMem_0_5_7 : _GEN_5626; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5628 = _GEN_9835 & _GEN_18226 ? CacheMem_0_6_7 : _GEN_5627; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5629 = _GEN_9835 & _GEN_18228 ? CacheMem_0_7_7 : _GEN_5628; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5630 = _GEN_10087 & _GEN_18230 ? CacheMem_1_0_7 : _GEN_5629; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5631 = _GEN_10087 & _GEN_18216 ? CacheMem_1_1_7 : _GEN_5630; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5632 = _GEN_10087 & _GEN_18218 ? CacheMem_1_2_7 : _GEN_5631; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5633 = _GEN_10087 & _GEN_18220 ? CacheMem_1_3_7 : _GEN_5632; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5634 = _GEN_10087 & _GEN_18222 ? CacheMem_1_4_7 : _GEN_5633; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5635 = _GEN_10087 & _GEN_18224 ? CacheMem_1_5_7 : _GEN_5634; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5636 = _GEN_10087 & _GEN_18226 ? CacheMem_1_6_7 : _GEN_5635; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5637 = _GEN_10087 & _GEN_18228 ? CacheMem_1_7_7 : _GEN_5636; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5638 = _GEN_10343 & _GEN_18230 ? CacheMem_2_0_7 : _GEN_5637; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5639 = _GEN_10343 & _GEN_18216 ? CacheMem_2_1_7 : _GEN_5638; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5640 = _GEN_10343 & _GEN_18218 ? CacheMem_2_2_7 : _GEN_5639; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5641 = _GEN_10343 & _GEN_18220 ? CacheMem_2_3_7 : _GEN_5640; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5642 = _GEN_10343 & _GEN_18222 ? CacheMem_2_4_7 : _GEN_5641; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5643 = _GEN_10343 & _GEN_18224 ? CacheMem_2_5_7 : _GEN_5642; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5644 = _GEN_10343 & _GEN_18226 ? CacheMem_2_6_7 : _GEN_5643; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5645 = _GEN_10343 & _GEN_18228 ? CacheMem_2_7_7 : _GEN_5644; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5646 = _GEN_10599 & _GEN_18230 ? CacheMem_3_0_7 : _GEN_5645; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5647 = _GEN_10599 & _GEN_18216 ? CacheMem_3_1_7 : _GEN_5646; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5648 = _GEN_10599 & _GEN_18218 ? CacheMem_3_2_7 : _GEN_5647; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5649 = _GEN_10599 & _GEN_18220 ? CacheMem_3_3_7 : _GEN_5648; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5650 = _GEN_10599 & _GEN_18222 ? CacheMem_3_4_7 : _GEN_5649; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5651 = _GEN_10599 & _GEN_18224 ? CacheMem_3_5_7 : _GEN_5650; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5652 = _GEN_10599 & _GEN_18226 ? CacheMem_3_6_7 : _GEN_5651; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5653 = _GEN_10599 & _GEN_18228 ? CacheMem_3_7_7 : _GEN_5652; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5654 = _GEN_10855 & _GEN_18230 ? CacheMem_4_0_7 : _GEN_5653; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5655 = _GEN_10855 & _GEN_18216 ? CacheMem_4_1_7 : _GEN_5654; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5656 = _GEN_10855 & _GEN_18218 ? CacheMem_4_2_7 : _GEN_5655; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5657 = _GEN_10855 & _GEN_18220 ? CacheMem_4_3_7 : _GEN_5656; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5658 = _GEN_10855 & _GEN_18222 ? CacheMem_4_4_7 : _GEN_5657; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5659 = _GEN_10855 & _GEN_18224 ? CacheMem_4_5_7 : _GEN_5658; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5660 = _GEN_10855 & _GEN_18226 ? CacheMem_4_6_7 : _GEN_5659; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5661 = _GEN_10855 & _GEN_18228 ? CacheMem_4_7_7 : _GEN_5660; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5662 = _GEN_11111 & _GEN_18230 ? CacheMem_5_0_7 : _GEN_5661; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5663 = _GEN_11111 & _GEN_18216 ? CacheMem_5_1_7 : _GEN_5662; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5664 = _GEN_11111 & _GEN_18218 ? CacheMem_5_2_7 : _GEN_5663; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5665 = _GEN_11111 & _GEN_18220 ? CacheMem_5_3_7 : _GEN_5664; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5666 = _GEN_11111 & _GEN_18222 ? CacheMem_5_4_7 : _GEN_5665; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5667 = _GEN_11111 & _GEN_18224 ? CacheMem_5_5_7 : _GEN_5666; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5668 = _GEN_11111 & _GEN_18226 ? CacheMem_5_6_7 : _GEN_5667; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5669 = _GEN_11111 & _GEN_18228 ? CacheMem_5_7_7 : _GEN_5668; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5670 = _GEN_11367 & _GEN_18230 ? CacheMem_6_0_7 : _GEN_5669; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5671 = _GEN_11367 & _GEN_18216 ? CacheMem_6_1_7 : _GEN_5670; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5672 = _GEN_11367 & _GEN_18218 ? CacheMem_6_2_7 : _GEN_5671; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5673 = _GEN_11367 & _GEN_18220 ? CacheMem_6_3_7 : _GEN_5672; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5674 = _GEN_11367 & _GEN_18222 ? CacheMem_6_4_7 : _GEN_5673; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5675 = _GEN_11367 & _GEN_18224 ? CacheMem_6_5_7 : _GEN_5674; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5676 = _GEN_11367 & _GEN_18226 ? CacheMem_6_6_7 : _GEN_5675; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5677 = _GEN_11367 & _GEN_18228 ? CacheMem_6_7_7 : _GEN_5676; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5678 = _GEN_11623 & _GEN_18230 ? CacheMem_7_0_7 : _GEN_5677; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5679 = _GEN_11623 & _GEN_18216 ? CacheMem_7_1_7 : _GEN_5678; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5680 = _GEN_11623 & _GEN_18218 ? CacheMem_7_2_7 : _GEN_5679; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5681 = _GEN_11623 & _GEN_18220 ? CacheMem_7_3_7 : _GEN_5680; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5682 = _GEN_11623 & _GEN_18222 ? CacheMem_7_4_7 : _GEN_5681; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5683 = _GEN_11623 & _GEN_18224 ? CacheMem_7_5_7 : _GEN_5682; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5684 = _GEN_11623 & _GEN_18226 ? CacheMem_7_6_7 : _GEN_5683; // @[Cache.scala 153:{25,25}]
  wire [31:0] _GEN_5685 = _GEN_11623 & _GEN_18228 ? CacheMem_7_7_7 : _GEN_5684; // @[Cache.scala 153:{25,25}]
  wire [1:0] _GEN_5686 = _GEN_5045 & _GEN_5109 ? 2'h1 : 2'h2; // @[Cache.scala 150:103 151:24 155:24]
  wire [8:0] _GEN_5687 = _GEN_5045 & _GEN_5109 ? _mem_wr_addr_T : mem_wr_addr; // @[Cache.scala 150:103 152:25 73:28]
  wire [31:0] _GEN_5688 = _GEN_5045 & _GEN_5109 ? _GEN_5237 : mem_wr_line_0; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5689 = _GEN_5045 & _GEN_5109 ? _GEN_5301 : mem_wr_line_1; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5690 = _GEN_5045 & _GEN_5109 ? _GEN_5365 : mem_wr_line_2; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5691 = _GEN_5045 & _GEN_5109 ? _GEN_5429 : mem_wr_line_3; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5692 = _GEN_5045 & _GEN_5109 ? _GEN_5493 : mem_wr_line_4; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5693 = _GEN_5045 & _GEN_5109 ? _GEN_5557 : mem_wr_line_5; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5694 = _GEN_5045 & _GEN_5109 ? _GEN_5621 : mem_wr_line_6; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5695 = _GEN_5045 & _GEN_5109 ? _GEN_5685 : mem_wr_line_7; // @[Cache.scala 150:103 153:25 124:28]
  wire [31:0] _GEN_5708 = cache_Hit ? _GEN_4404 : 32'h0; // @[Cache.scala 128:22]
  wire [1:0] _GEN_6298 = io_cacheAXI_gnt ? 2'h3 : cacheState; // @[Cache.scala 168:39 169:20 96:27]
  wire  _GEN_19601 = 3'h0 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6299 = 3'h0 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_0_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6300 = 3'h0 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_0_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6301 = 3'h0 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_0_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6302 = 3'h0 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_0_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6303 = 3'h0 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_0_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6304 = 3'h0 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_0_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6305 = 3'h0 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_0_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6306 = 3'h0 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_0_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19617 = 3'h1 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6307 = 3'h1 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_1_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6308 = 3'h1 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_1_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6309 = 3'h1 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_1_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6310 = 3'h1 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_1_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6311 = 3'h1 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_1_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6312 = 3'h1 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_1_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6313 = 3'h1 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_1_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6314 = 3'h1 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_1_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19633 = 3'h2 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6315 = 3'h2 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_2_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6316 = 3'h2 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_2_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6317 = 3'h2 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_2_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6318 = 3'h2 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_2_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6319 = 3'h2 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_2_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6320 = 3'h2 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_2_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6321 = 3'h2 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_2_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6322 = 3'h2 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_2_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19649 = 3'h3 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6323 = 3'h3 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_3_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6324 = 3'h3 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_3_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6325 = 3'h3 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_3_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6326 = 3'h3 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_3_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6327 = 3'h3 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_3_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6328 = 3'h3 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_3_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6329 = 3'h3 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_3_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6330 = 3'h3 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_3_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19665 = 3'h4 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6331 = 3'h4 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_4_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6332 = 3'h4 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_4_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6333 = 3'h4 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_4_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6334 = 3'h4 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_4_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6335 = 3'h4 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_4_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6336 = 3'h4 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_4_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6337 = 3'h4 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_4_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6338 = 3'h4 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_4_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19681 = 3'h5 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6339 = 3'h5 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_5_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6340 = 3'h5 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_5_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6341 = 3'h5 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_5_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6342 = 3'h5 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_5_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6343 = 3'h5 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_5_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6344 = 3'h5 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_5_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6345 = 3'h5 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_5_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6346 = 3'h5 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_5_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19697 = 3'h6 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6347 = 3'h6 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_6_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6348 = 3'h6 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_6_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6349 = 3'h6 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_6_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6350 = 3'h6 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_6_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6351 = 3'h6 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_6_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6352 = 3'h6 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_6_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6353 = 3'h6 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_6_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6354 = 3'h6 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_6_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_19713 = 3'h7 == mem_rd_set_addr; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6355 = 3'h7 == mem_rd_set_addr & _GEN_18230 ? mem_rd_tag_addr : cache_tags_7_0; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6356 = 3'h7 == mem_rd_set_addr & _GEN_18216 ? mem_rd_tag_addr : cache_tags_7_1; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6357 = 3'h7 == mem_rd_set_addr & _GEN_18218 ? mem_rd_tag_addr : cache_tags_7_2; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6358 = 3'h7 == mem_rd_set_addr & _GEN_18220 ? mem_rd_tag_addr : cache_tags_7_3; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6359 = 3'h7 == mem_rd_set_addr & _GEN_18222 ? mem_rd_tag_addr : cache_tags_7_4; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6360 = 3'h7 == mem_rd_set_addr & _GEN_18224 ? mem_rd_tag_addr : cache_tags_7_5; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6361 = 3'h7 == mem_rd_set_addr & _GEN_18226 ? mem_rd_tag_addr : cache_tags_7_6; // @[Cache.scala 174:{50,50} 56:27]
  wire [5:0] _GEN_6362 = 3'h7 == mem_rd_set_addr & _GEN_18228 ? mem_rd_tag_addr : cache_tags_7_7; // @[Cache.scala 174:{50,50} 56:27]
  wire  _GEN_6363 = _GEN_19601 & _GEN_18230 | valid_0_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6364 = _GEN_19601 & _GEN_18216 | valid_0_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6365 = _GEN_19601 & _GEN_18218 | valid_0_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6366 = _GEN_19601 & _GEN_18220 | valid_0_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6367 = _GEN_19601 & _GEN_18222 | valid_0_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6368 = _GEN_19601 & _GEN_18224 | valid_0_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6369 = _GEN_19601 & _GEN_18226 | valid_0_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6370 = _GEN_19601 & _GEN_18228 | valid_0_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6371 = _GEN_19617 & _GEN_18230 | valid_1_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6372 = _GEN_19617 & _GEN_18216 | valid_1_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6373 = _GEN_19617 & _GEN_18218 | valid_1_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6374 = _GEN_19617 & _GEN_18220 | valid_1_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6375 = _GEN_19617 & _GEN_18222 | valid_1_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6376 = _GEN_19617 & _GEN_18224 | valid_1_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6377 = _GEN_19617 & _GEN_18226 | valid_1_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6378 = _GEN_19617 & _GEN_18228 | valid_1_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6379 = _GEN_19633 & _GEN_18230 | valid_2_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6380 = _GEN_19633 & _GEN_18216 | valid_2_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6381 = _GEN_19633 & _GEN_18218 | valid_2_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6382 = _GEN_19633 & _GEN_18220 | valid_2_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6383 = _GEN_19633 & _GEN_18222 | valid_2_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6384 = _GEN_19633 & _GEN_18224 | valid_2_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6385 = _GEN_19633 & _GEN_18226 | valid_2_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6386 = _GEN_19633 & _GEN_18228 | valid_2_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6387 = _GEN_19649 & _GEN_18230 | valid_3_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6388 = _GEN_19649 & _GEN_18216 | valid_3_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6389 = _GEN_19649 & _GEN_18218 | valid_3_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6390 = _GEN_19649 & _GEN_18220 | valid_3_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6391 = _GEN_19649 & _GEN_18222 | valid_3_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6392 = _GEN_19649 & _GEN_18224 | valid_3_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6393 = _GEN_19649 & _GEN_18226 | valid_3_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6394 = _GEN_19649 & _GEN_18228 | valid_3_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6395 = _GEN_19665 & _GEN_18230 | valid_4_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6396 = _GEN_19665 & _GEN_18216 | valid_4_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6397 = _GEN_19665 & _GEN_18218 | valid_4_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6398 = _GEN_19665 & _GEN_18220 | valid_4_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6399 = _GEN_19665 & _GEN_18222 | valid_4_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6400 = _GEN_19665 & _GEN_18224 | valid_4_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6401 = _GEN_19665 & _GEN_18226 | valid_4_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6402 = _GEN_19665 & _GEN_18228 | valid_4_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6403 = _GEN_19681 & _GEN_18230 | valid_5_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6404 = _GEN_19681 & _GEN_18216 | valid_5_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6405 = _GEN_19681 & _GEN_18218 | valid_5_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6406 = _GEN_19681 & _GEN_18220 | valid_5_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6407 = _GEN_19681 & _GEN_18222 | valid_5_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6408 = _GEN_19681 & _GEN_18224 | valid_5_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6409 = _GEN_19681 & _GEN_18226 | valid_5_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6410 = _GEN_19681 & _GEN_18228 | valid_5_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6411 = _GEN_19697 & _GEN_18230 | valid_6_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6412 = _GEN_19697 & _GEN_18216 | valid_6_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6413 = _GEN_19697 & _GEN_18218 | valid_6_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6414 = _GEN_19697 & _GEN_18220 | valid_6_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6415 = _GEN_19697 & _GEN_18222 | valid_6_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6416 = _GEN_19697 & _GEN_18224 | valid_6_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6417 = _GEN_19697 & _GEN_18226 | valid_6_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6418 = _GEN_19697 & _GEN_18228 | valid_6_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6419 = _GEN_19713 & _GEN_18230 | valid_7_0; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6420 = _GEN_19713 & _GEN_18216 | valid_7_1; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6421 = _GEN_19713 & _GEN_18218 | valid_7_2; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6422 = _GEN_19713 & _GEN_18220 | valid_7_3; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6423 = _GEN_19713 & _GEN_18222 | valid_7_4; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6424 = _GEN_19713 & _GEN_18224 | valid_7_5; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6425 = _GEN_19713 & _GEN_18226 | valid_7_6; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6426 = _GEN_19713 & _GEN_18228 | valid_7_7; // @[Cache.scala 175:{45,45} 57:22]
  wire  _GEN_6427 = _GEN_19601 & _GEN_18230 ? 1'h0 : dirty_0_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6428 = _GEN_19601 & _GEN_18216 ? 1'h0 : dirty_0_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6429 = _GEN_19601 & _GEN_18218 ? 1'h0 : dirty_0_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6430 = _GEN_19601 & _GEN_18220 ? 1'h0 : dirty_0_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6431 = _GEN_19601 & _GEN_18222 ? 1'h0 : dirty_0_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6432 = _GEN_19601 & _GEN_18224 ? 1'h0 : dirty_0_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6433 = _GEN_19601 & _GEN_18226 ? 1'h0 : dirty_0_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6434 = _GEN_19601 & _GEN_18228 ? 1'h0 : dirty_0_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6435 = _GEN_19617 & _GEN_18230 ? 1'h0 : dirty_1_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6436 = _GEN_19617 & _GEN_18216 ? 1'h0 : dirty_1_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6437 = _GEN_19617 & _GEN_18218 ? 1'h0 : dirty_1_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6438 = _GEN_19617 & _GEN_18220 ? 1'h0 : dirty_1_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6439 = _GEN_19617 & _GEN_18222 ? 1'h0 : dirty_1_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6440 = _GEN_19617 & _GEN_18224 ? 1'h0 : dirty_1_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6441 = _GEN_19617 & _GEN_18226 ? 1'h0 : dirty_1_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6442 = _GEN_19617 & _GEN_18228 ? 1'h0 : dirty_1_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6443 = _GEN_19633 & _GEN_18230 ? 1'h0 : dirty_2_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6444 = _GEN_19633 & _GEN_18216 ? 1'h0 : dirty_2_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6445 = _GEN_19633 & _GEN_18218 ? 1'h0 : dirty_2_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6446 = _GEN_19633 & _GEN_18220 ? 1'h0 : dirty_2_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6447 = _GEN_19633 & _GEN_18222 ? 1'h0 : dirty_2_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6448 = _GEN_19633 & _GEN_18224 ? 1'h0 : dirty_2_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6449 = _GEN_19633 & _GEN_18226 ? 1'h0 : dirty_2_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6450 = _GEN_19633 & _GEN_18228 ? 1'h0 : dirty_2_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6451 = _GEN_19649 & _GEN_18230 ? 1'h0 : dirty_3_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6452 = _GEN_19649 & _GEN_18216 ? 1'h0 : dirty_3_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6453 = _GEN_19649 & _GEN_18218 ? 1'h0 : dirty_3_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6454 = _GEN_19649 & _GEN_18220 ? 1'h0 : dirty_3_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6455 = _GEN_19649 & _GEN_18222 ? 1'h0 : dirty_3_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6456 = _GEN_19649 & _GEN_18224 ? 1'h0 : dirty_3_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6457 = _GEN_19649 & _GEN_18226 ? 1'h0 : dirty_3_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6458 = _GEN_19649 & _GEN_18228 ? 1'h0 : dirty_3_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6459 = _GEN_19665 & _GEN_18230 ? 1'h0 : dirty_4_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6460 = _GEN_19665 & _GEN_18216 ? 1'h0 : dirty_4_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6461 = _GEN_19665 & _GEN_18218 ? 1'h0 : dirty_4_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6462 = _GEN_19665 & _GEN_18220 ? 1'h0 : dirty_4_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6463 = _GEN_19665 & _GEN_18222 ? 1'h0 : dirty_4_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6464 = _GEN_19665 & _GEN_18224 ? 1'h0 : dirty_4_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6465 = _GEN_19665 & _GEN_18226 ? 1'h0 : dirty_4_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6466 = _GEN_19665 & _GEN_18228 ? 1'h0 : dirty_4_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6467 = _GEN_19681 & _GEN_18230 ? 1'h0 : dirty_5_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6468 = _GEN_19681 & _GEN_18216 ? 1'h0 : dirty_5_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6469 = _GEN_19681 & _GEN_18218 ? 1'h0 : dirty_5_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6470 = _GEN_19681 & _GEN_18220 ? 1'h0 : dirty_5_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6471 = _GEN_19681 & _GEN_18222 ? 1'h0 : dirty_5_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6472 = _GEN_19681 & _GEN_18224 ? 1'h0 : dirty_5_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6473 = _GEN_19681 & _GEN_18226 ? 1'h0 : dirty_5_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6474 = _GEN_19681 & _GEN_18228 ? 1'h0 : dirty_5_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6475 = _GEN_19697 & _GEN_18230 ? 1'h0 : dirty_6_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6476 = _GEN_19697 & _GEN_18216 ? 1'h0 : dirty_6_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6477 = _GEN_19697 & _GEN_18218 ? 1'h0 : dirty_6_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6478 = _GEN_19697 & _GEN_18220 ? 1'h0 : dirty_6_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6479 = _GEN_19697 & _GEN_18222 ? 1'h0 : dirty_6_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6480 = _GEN_19697 & _GEN_18224 ? 1'h0 : dirty_6_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6481 = _GEN_19697 & _GEN_18226 ? 1'h0 : dirty_6_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6482 = _GEN_19697 & _GEN_18228 ? 1'h0 : dirty_6_7; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6483 = _GEN_19713 & _GEN_18230 ? 1'h0 : dirty_7_0; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6484 = _GEN_19713 & _GEN_18216 ? 1'h0 : dirty_7_1; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6485 = _GEN_19713 & _GEN_18218 ? 1'h0 : dirty_7_2; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6486 = _GEN_19713 & _GEN_18220 ? 1'h0 : dirty_7_3; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6487 = _GEN_19713 & _GEN_18222 ? 1'h0 : dirty_7_4; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6488 = _GEN_19713 & _GEN_18224 ? 1'h0 : dirty_7_5; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6489 = _GEN_19713 & _GEN_18226 ? 1'h0 : dirty_7_6; // @[Cache.scala 176:{45,45} 58:22]
  wire  _GEN_6490 = _GEN_19713 & _GEN_18228 ? 1'h0 : dirty_7_7; // @[Cache.scala 176:{45,45} 58:22]
  wire [31:0] _GEN_6491 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_0_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6492 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_0_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6493 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_0_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6494 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_0_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6495 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_0_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6496 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_0_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6497 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_0_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6498 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_0_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6499 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_1_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6500 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_1_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6501 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_1_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6502 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_1_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6503 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_1_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6504 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_1_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6505 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_1_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6506 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_1_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6507 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_2_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6508 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_2_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6509 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_2_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6510 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_2_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6511 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_2_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6512 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_2_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6513 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_2_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6514 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_2_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6515 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_3_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6516 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_3_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6517 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_3_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6518 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_3_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6519 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_3_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6520 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_3_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6521 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_3_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6522 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_3_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6523 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_4_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6524 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_4_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6525 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_4_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6526 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_4_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6527 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_4_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6528 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_4_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6529 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_4_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6530 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_4_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6531 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_5_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6532 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_5_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6533 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_5_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6534 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_5_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6535 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_5_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6536 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_5_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6537 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_5_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6538 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_5_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6539 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_6_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6540 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_6_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6541 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_6_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6542 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_6_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6543 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_6_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6544 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_6_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6545 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_6_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6546 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_6_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6547 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_0 : CacheMem_7_0_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6548 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_0 : CacheMem_7_1_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6549 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_0 : CacheMem_7_2_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6550 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_0 : CacheMem_7_3_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6551 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_0 : CacheMem_7_4_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6552 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_0 : CacheMem_7_5_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6553 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_0 : CacheMem_7_6_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6554 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_0 : CacheMem_7_7_0; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6555 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_0_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6556 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_0_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6557 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_0_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6558 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_0_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6559 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_0_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6560 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_0_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6561 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_0_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6562 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_0_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6563 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_1_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6564 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_1_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6565 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_1_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6566 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_1_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6567 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_1_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6568 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_1_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6569 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_1_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6570 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_1_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6571 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_2_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6572 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_2_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6573 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_2_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6574 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_2_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6575 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_2_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6576 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_2_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6577 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_2_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6578 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_2_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6579 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_3_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6580 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_3_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6581 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_3_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6582 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_3_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6583 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_3_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6584 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_3_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6585 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_3_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6586 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_3_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6587 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_4_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6588 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_4_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6589 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_4_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6590 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_4_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6591 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_4_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6592 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_4_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6593 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_4_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6594 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_4_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6595 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_5_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6596 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_5_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6597 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_5_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6598 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_5_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6599 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_5_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6600 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_5_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6601 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_5_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6602 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_5_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6603 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_6_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6604 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_6_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6605 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_6_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6606 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_6_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6607 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_6_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6608 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_6_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6609 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_6_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6610 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_6_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6611 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_1 : CacheMem_7_0_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6612 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_1 : CacheMem_7_1_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6613 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_1 : CacheMem_7_2_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6614 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_1 : CacheMem_7_3_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6615 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_1 : CacheMem_7_4_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6616 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_1 : CacheMem_7_5_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6617 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_1 : CacheMem_7_6_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6618 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_1 : CacheMem_7_7_1; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6619 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_0_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6620 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_0_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6621 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_0_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6622 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_0_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6623 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_0_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6624 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_0_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6625 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_0_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6626 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_0_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6627 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_1_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6628 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_1_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6629 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_1_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6630 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_1_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6631 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_1_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6632 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_1_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6633 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_1_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6634 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_1_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6635 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_2_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6636 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_2_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6637 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_2_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6638 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_2_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6639 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_2_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6640 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_2_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6641 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_2_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6642 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_2_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6643 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_3_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6644 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_3_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6645 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_3_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6646 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_3_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6647 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_3_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6648 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_3_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6649 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_3_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6650 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_3_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6651 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_4_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6652 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_4_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6653 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_4_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6654 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_4_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6655 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_4_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6656 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_4_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6657 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_4_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6658 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_4_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6659 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_5_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6660 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_5_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6661 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_5_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6662 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_5_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6663 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_5_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6664 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_5_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6665 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_5_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6666 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_5_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6667 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_6_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6668 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_6_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6669 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_6_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6670 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_6_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6671 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_6_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6672 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_6_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6673 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_6_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6674 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_6_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6675 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_2 : CacheMem_7_0_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6676 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_2 : CacheMem_7_1_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6677 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_2 : CacheMem_7_2_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6678 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_2 : CacheMem_7_3_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6679 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_2 : CacheMem_7_4_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6680 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_2 : CacheMem_7_5_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6681 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_2 : CacheMem_7_6_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6682 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_2 : CacheMem_7_7_2; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6683 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_0_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6684 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_0_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6685 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_0_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6686 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_0_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6687 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_0_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6688 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_0_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6689 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_0_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6690 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_0_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6691 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_1_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6692 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_1_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6693 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_1_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6694 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_1_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6695 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_1_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6696 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_1_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6697 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_1_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6698 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_1_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6699 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_2_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6700 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_2_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6701 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_2_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6702 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_2_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6703 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_2_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6704 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_2_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6705 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_2_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6706 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_2_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6707 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_3_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6708 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_3_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6709 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_3_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6710 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_3_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6711 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_3_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6712 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_3_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6713 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_3_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6714 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_3_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6715 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_4_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6716 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_4_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6717 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_4_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6718 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_4_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6719 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_4_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6720 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_4_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6721 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_4_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6722 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_4_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6723 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_5_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6724 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_5_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6725 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_5_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6726 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_5_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6727 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_5_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6728 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_5_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6729 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_5_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6730 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_5_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6731 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_6_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6732 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_6_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6733 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_6_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6734 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_6_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6735 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_6_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6736 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_6_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6737 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_6_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6738 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_6_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6739 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_3 : CacheMem_7_0_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6740 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_3 : CacheMem_7_1_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6741 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_3 : CacheMem_7_2_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6742 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_3 : CacheMem_7_3_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6743 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_3 : CacheMem_7_4_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6744 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_3 : CacheMem_7_5_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6745 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_3 : CacheMem_7_6_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6746 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_3 : CacheMem_7_7_3; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6747 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_0_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6748 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_0_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6749 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_0_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6750 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_0_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6751 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_0_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6752 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_0_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6753 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_0_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6754 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_0_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6755 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_1_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6756 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_1_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6757 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_1_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6758 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_1_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6759 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_1_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6760 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_1_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6761 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_1_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6762 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_1_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6763 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_2_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6764 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_2_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6765 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_2_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6766 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_2_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6767 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_2_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6768 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_2_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6769 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_2_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6770 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_2_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6771 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_3_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6772 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_3_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6773 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_3_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6774 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_3_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6775 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_3_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6776 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_3_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6777 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_3_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6778 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_3_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6779 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_4_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6780 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_4_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6781 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_4_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6782 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_4_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6783 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_4_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6784 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_4_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6785 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_4_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6786 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_4_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6787 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_5_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6788 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_5_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6789 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_5_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6790 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_5_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6791 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_5_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6792 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_5_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6793 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_5_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6794 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_5_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6795 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_6_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6796 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_6_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6797 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_6_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6798 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_6_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6799 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_6_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6800 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_6_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6801 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_6_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6802 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_6_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6803 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_4 : CacheMem_7_0_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6804 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_4 : CacheMem_7_1_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6805 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_4 : CacheMem_7_2_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6806 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_4 : CacheMem_7_3_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6807 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_4 : CacheMem_7_4_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6808 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_4 : CacheMem_7_5_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6809 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_4 : CacheMem_7_6_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6810 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_4 : CacheMem_7_7_4; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6811 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_0_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6812 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_0_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6813 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_0_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6814 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_0_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6815 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_0_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6816 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_0_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6817 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_0_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6818 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_0_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6819 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_1_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6820 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_1_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6821 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_1_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6822 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_1_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6823 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_1_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6824 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_1_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6825 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_1_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6826 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_1_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6827 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_2_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6828 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_2_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6829 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_2_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6830 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_2_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6831 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_2_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6832 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_2_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6833 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_2_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6834 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_2_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6835 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_3_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6836 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_3_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6837 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_3_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6838 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_3_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6839 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_3_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6840 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_3_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6841 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_3_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6842 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_3_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6843 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_4_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6844 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_4_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6845 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_4_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6846 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_4_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6847 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_4_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6848 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_4_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6849 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_4_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6850 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_4_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6851 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_5_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6852 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_5_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6853 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_5_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6854 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_5_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6855 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_5_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6856 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_5_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6857 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_5_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6858 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_5_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6859 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_6_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6860 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_6_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6861 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_6_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6862 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_6_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6863 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_6_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6864 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_6_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6865 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_6_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6866 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_6_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6867 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_5 : CacheMem_7_0_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6868 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_5 : CacheMem_7_1_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6869 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_5 : CacheMem_7_2_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6870 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_5 : CacheMem_7_3_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6871 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_5 : CacheMem_7_4_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6872 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_5 : CacheMem_7_5_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6873 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_5 : CacheMem_7_6_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6874 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_5 : CacheMem_7_7_5; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6875 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_0_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6876 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_0_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6877 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_0_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6878 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_0_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6879 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_0_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6880 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_0_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6881 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_0_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6882 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_0_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6883 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_1_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6884 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_1_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6885 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_1_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6886 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_1_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6887 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_1_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6888 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_1_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6889 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_1_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6890 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_1_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6891 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_2_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6892 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_2_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6893 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_2_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6894 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_2_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6895 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_2_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6896 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_2_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6897 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_2_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6898 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_2_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6899 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_3_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6900 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_3_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6901 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_3_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6902 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_3_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6903 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_3_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6904 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_3_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6905 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_3_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6906 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_3_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6907 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_4_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6908 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_4_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6909 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_4_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6910 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_4_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6911 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_4_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6912 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_4_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6913 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_4_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6914 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_4_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6915 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_5_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6916 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_5_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6917 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_5_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6918 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_5_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6919 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_5_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6920 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_5_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6921 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_5_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6922 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_5_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6923 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_6_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6924 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_6_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6925 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_6_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6926 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_6_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6927 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_6_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6928 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_6_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6929 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_6_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6930 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_6_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6931 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_6 : CacheMem_7_0_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6932 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_6 : CacheMem_7_1_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6933 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_6 : CacheMem_7_2_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6934 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_6 : CacheMem_7_3_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6935 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_6 : CacheMem_7_4_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6936 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_6 : CacheMem_7_5_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6937 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_6 : CacheMem_7_6_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6938 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_6 : CacheMem_7_7_6; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6939 = _GEN_19601 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_0_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6940 = _GEN_19601 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_0_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6941 = _GEN_19601 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_0_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6942 = _GEN_19601 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_0_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6943 = _GEN_19601 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_0_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6944 = _GEN_19601 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_0_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6945 = _GEN_19601 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_0_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6946 = _GEN_19601 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_0_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6947 = _GEN_19617 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_1_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6948 = _GEN_19617 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_1_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6949 = _GEN_19617 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_1_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6950 = _GEN_19617 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_1_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6951 = _GEN_19617 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_1_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6952 = _GEN_19617 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_1_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6953 = _GEN_19617 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_1_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6954 = _GEN_19617 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_1_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6955 = _GEN_19633 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_2_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6956 = _GEN_19633 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_2_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6957 = _GEN_19633 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_2_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6958 = _GEN_19633 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_2_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6959 = _GEN_19633 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_2_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6960 = _GEN_19633 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_2_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6961 = _GEN_19633 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_2_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6962 = _GEN_19633 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_2_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6963 = _GEN_19649 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_3_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6964 = _GEN_19649 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_3_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6965 = _GEN_19649 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_3_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6966 = _GEN_19649 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_3_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6967 = _GEN_19649 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_3_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6968 = _GEN_19649 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_3_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6969 = _GEN_19649 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_3_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6970 = _GEN_19649 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_3_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6971 = _GEN_19665 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_4_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6972 = _GEN_19665 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_4_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6973 = _GEN_19665 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_4_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6974 = _GEN_19665 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_4_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6975 = _GEN_19665 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_4_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6976 = _GEN_19665 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_4_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6977 = _GEN_19665 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_4_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6978 = _GEN_19665 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_4_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6979 = _GEN_19681 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_5_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6980 = _GEN_19681 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_5_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6981 = _GEN_19681 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_5_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6982 = _GEN_19681 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_5_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6983 = _GEN_19681 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_5_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6984 = _GEN_19681 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_5_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6985 = _GEN_19681 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_5_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6986 = _GEN_19681 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_5_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6987 = _GEN_19697 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_6_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6988 = _GEN_19697 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_6_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6989 = _GEN_19697 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_6_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6990 = _GEN_19697 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_6_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6991 = _GEN_19697 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_6_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6992 = _GEN_19697 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_6_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6993 = _GEN_19697 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_6_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6994 = _GEN_19697 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_6_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6995 = _GEN_19713 & _GEN_18230 ? io_mem_rd_line_7 : CacheMem_7_0_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6996 = _GEN_19713 & _GEN_18216 ? io_mem_rd_line_7 : CacheMem_7_1_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6997 = _GEN_19713 & _GEN_18218 ? io_mem_rd_line_7 : CacheMem_7_2_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6998 = _GEN_19713 & _GEN_18220 ? io_mem_rd_line_7 : CacheMem_7_3_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_6999 = _GEN_19713 & _GEN_18222 ? io_mem_rd_line_7 : CacheMem_7_4_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_7000 = _GEN_19713 & _GEN_18224 ? io_mem_rd_line_7 : CacheMem_7_5_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_7001 = _GEN_19713 & _GEN_18226 ? io_mem_rd_line_7 : CacheMem_7_6_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [31:0] _GEN_7002 = _GEN_19713 & _GEN_18228 ? io_mem_rd_line_7 : CacheMem_7_7_7; // @[Cache.scala 178:{55,55} 53:25]
  wire [1:0] _GEN_7003 = _T_30 ? 2'h0 : cacheState; // @[Cache.scala 126:21 173:18 96:27]
  wire [5:0] _GEN_7004 = _T_30 ? _GEN_6299 : cache_tags_0_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7005 = _T_30 ? _GEN_6300 : cache_tags_0_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7006 = _T_30 ? _GEN_6301 : cache_tags_0_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7007 = _T_30 ? _GEN_6302 : cache_tags_0_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7008 = _T_30 ? _GEN_6303 : cache_tags_0_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7009 = _T_30 ? _GEN_6304 : cache_tags_0_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7010 = _T_30 ? _GEN_6305 : cache_tags_0_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7011 = _T_30 ? _GEN_6306 : cache_tags_0_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7012 = _T_30 ? _GEN_6307 : cache_tags_1_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7013 = _T_30 ? _GEN_6308 : cache_tags_1_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7014 = _T_30 ? _GEN_6309 : cache_tags_1_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7015 = _T_30 ? _GEN_6310 : cache_tags_1_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7016 = _T_30 ? _GEN_6311 : cache_tags_1_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7017 = _T_30 ? _GEN_6312 : cache_tags_1_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7018 = _T_30 ? _GEN_6313 : cache_tags_1_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7019 = _T_30 ? _GEN_6314 : cache_tags_1_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7020 = _T_30 ? _GEN_6315 : cache_tags_2_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7021 = _T_30 ? _GEN_6316 : cache_tags_2_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7022 = _T_30 ? _GEN_6317 : cache_tags_2_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7023 = _T_30 ? _GEN_6318 : cache_tags_2_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7024 = _T_30 ? _GEN_6319 : cache_tags_2_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7025 = _T_30 ? _GEN_6320 : cache_tags_2_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7026 = _T_30 ? _GEN_6321 : cache_tags_2_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7027 = _T_30 ? _GEN_6322 : cache_tags_2_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7028 = _T_30 ? _GEN_6323 : cache_tags_3_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7029 = _T_30 ? _GEN_6324 : cache_tags_3_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7030 = _T_30 ? _GEN_6325 : cache_tags_3_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7031 = _T_30 ? _GEN_6326 : cache_tags_3_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7032 = _T_30 ? _GEN_6327 : cache_tags_3_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7033 = _T_30 ? _GEN_6328 : cache_tags_3_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7034 = _T_30 ? _GEN_6329 : cache_tags_3_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7035 = _T_30 ? _GEN_6330 : cache_tags_3_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7036 = _T_30 ? _GEN_6331 : cache_tags_4_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7037 = _T_30 ? _GEN_6332 : cache_tags_4_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7038 = _T_30 ? _GEN_6333 : cache_tags_4_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7039 = _T_30 ? _GEN_6334 : cache_tags_4_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7040 = _T_30 ? _GEN_6335 : cache_tags_4_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7041 = _T_30 ? _GEN_6336 : cache_tags_4_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7042 = _T_30 ? _GEN_6337 : cache_tags_4_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7043 = _T_30 ? _GEN_6338 : cache_tags_4_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7044 = _T_30 ? _GEN_6339 : cache_tags_5_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7045 = _T_30 ? _GEN_6340 : cache_tags_5_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7046 = _T_30 ? _GEN_6341 : cache_tags_5_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7047 = _T_30 ? _GEN_6342 : cache_tags_5_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7048 = _T_30 ? _GEN_6343 : cache_tags_5_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7049 = _T_30 ? _GEN_6344 : cache_tags_5_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7050 = _T_30 ? _GEN_6345 : cache_tags_5_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7051 = _T_30 ? _GEN_6346 : cache_tags_5_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7052 = _T_30 ? _GEN_6347 : cache_tags_6_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7053 = _T_30 ? _GEN_6348 : cache_tags_6_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7054 = _T_30 ? _GEN_6349 : cache_tags_6_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7055 = _T_30 ? _GEN_6350 : cache_tags_6_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7056 = _T_30 ? _GEN_6351 : cache_tags_6_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7057 = _T_30 ? _GEN_6352 : cache_tags_6_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7058 = _T_30 ? _GEN_6353 : cache_tags_6_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7059 = _T_30 ? _GEN_6354 : cache_tags_6_7; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7060 = _T_30 ? _GEN_6355 : cache_tags_7_0; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7061 = _T_30 ? _GEN_6356 : cache_tags_7_1; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7062 = _T_30 ? _GEN_6357 : cache_tags_7_2; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7063 = _T_30 ? _GEN_6358 : cache_tags_7_3; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7064 = _T_30 ? _GEN_6359 : cache_tags_7_4; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7065 = _T_30 ? _GEN_6360 : cache_tags_7_5; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7066 = _T_30 ? _GEN_6361 : cache_tags_7_6; // @[Cache.scala 126:21 56:27]
  wire [5:0] _GEN_7067 = _T_30 ? _GEN_6362 : cache_tags_7_7; // @[Cache.scala 126:21 56:27]
  wire  _GEN_7068 = _T_30 ? _GEN_6363 : valid_0_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7069 = _T_30 ? _GEN_6364 : valid_0_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7070 = _T_30 ? _GEN_6365 : valid_0_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7071 = _T_30 ? _GEN_6366 : valid_0_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7072 = _T_30 ? _GEN_6367 : valid_0_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7073 = _T_30 ? _GEN_6368 : valid_0_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7074 = _T_30 ? _GEN_6369 : valid_0_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7075 = _T_30 ? _GEN_6370 : valid_0_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7076 = _T_30 ? _GEN_6371 : valid_1_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7077 = _T_30 ? _GEN_6372 : valid_1_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7078 = _T_30 ? _GEN_6373 : valid_1_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7079 = _T_30 ? _GEN_6374 : valid_1_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7080 = _T_30 ? _GEN_6375 : valid_1_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7081 = _T_30 ? _GEN_6376 : valid_1_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7082 = _T_30 ? _GEN_6377 : valid_1_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7083 = _T_30 ? _GEN_6378 : valid_1_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7084 = _T_30 ? _GEN_6379 : valid_2_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7085 = _T_30 ? _GEN_6380 : valid_2_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7086 = _T_30 ? _GEN_6381 : valid_2_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7087 = _T_30 ? _GEN_6382 : valid_2_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7088 = _T_30 ? _GEN_6383 : valid_2_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7089 = _T_30 ? _GEN_6384 : valid_2_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7090 = _T_30 ? _GEN_6385 : valid_2_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7091 = _T_30 ? _GEN_6386 : valid_2_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7092 = _T_30 ? _GEN_6387 : valid_3_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7093 = _T_30 ? _GEN_6388 : valid_3_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7094 = _T_30 ? _GEN_6389 : valid_3_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7095 = _T_30 ? _GEN_6390 : valid_3_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7096 = _T_30 ? _GEN_6391 : valid_3_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7097 = _T_30 ? _GEN_6392 : valid_3_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7098 = _T_30 ? _GEN_6393 : valid_3_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7099 = _T_30 ? _GEN_6394 : valid_3_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7100 = _T_30 ? _GEN_6395 : valid_4_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7101 = _T_30 ? _GEN_6396 : valid_4_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7102 = _T_30 ? _GEN_6397 : valid_4_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7103 = _T_30 ? _GEN_6398 : valid_4_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7104 = _T_30 ? _GEN_6399 : valid_4_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7105 = _T_30 ? _GEN_6400 : valid_4_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7106 = _T_30 ? _GEN_6401 : valid_4_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7107 = _T_30 ? _GEN_6402 : valid_4_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7108 = _T_30 ? _GEN_6403 : valid_5_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7109 = _T_30 ? _GEN_6404 : valid_5_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7110 = _T_30 ? _GEN_6405 : valid_5_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7111 = _T_30 ? _GEN_6406 : valid_5_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7112 = _T_30 ? _GEN_6407 : valid_5_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7113 = _T_30 ? _GEN_6408 : valid_5_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7114 = _T_30 ? _GEN_6409 : valid_5_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7115 = _T_30 ? _GEN_6410 : valid_5_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7116 = _T_30 ? _GEN_6411 : valid_6_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7117 = _T_30 ? _GEN_6412 : valid_6_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7118 = _T_30 ? _GEN_6413 : valid_6_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7119 = _T_30 ? _GEN_6414 : valid_6_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7120 = _T_30 ? _GEN_6415 : valid_6_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7121 = _T_30 ? _GEN_6416 : valid_6_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7122 = _T_30 ? _GEN_6417 : valid_6_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7123 = _T_30 ? _GEN_6418 : valid_6_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7124 = _T_30 ? _GEN_6419 : valid_7_0; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7125 = _T_30 ? _GEN_6420 : valid_7_1; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7126 = _T_30 ? _GEN_6421 : valid_7_2; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7127 = _T_30 ? _GEN_6422 : valid_7_3; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7128 = _T_30 ? _GEN_6423 : valid_7_4; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7129 = _T_30 ? _GEN_6424 : valid_7_5; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7130 = _T_30 ? _GEN_6425 : valid_7_6; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7131 = _T_30 ? _GEN_6426 : valid_7_7; // @[Cache.scala 126:21 57:22]
  wire  _GEN_7132 = _T_30 ? _GEN_6427 : dirty_0_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7133 = _T_30 ? _GEN_6428 : dirty_0_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7134 = _T_30 ? _GEN_6429 : dirty_0_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7135 = _T_30 ? _GEN_6430 : dirty_0_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7136 = _T_30 ? _GEN_6431 : dirty_0_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7137 = _T_30 ? _GEN_6432 : dirty_0_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7138 = _T_30 ? _GEN_6433 : dirty_0_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7139 = _T_30 ? _GEN_6434 : dirty_0_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7140 = _T_30 ? _GEN_6435 : dirty_1_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7141 = _T_30 ? _GEN_6436 : dirty_1_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7142 = _T_30 ? _GEN_6437 : dirty_1_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7143 = _T_30 ? _GEN_6438 : dirty_1_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7144 = _T_30 ? _GEN_6439 : dirty_1_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7145 = _T_30 ? _GEN_6440 : dirty_1_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7146 = _T_30 ? _GEN_6441 : dirty_1_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7147 = _T_30 ? _GEN_6442 : dirty_1_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7148 = _T_30 ? _GEN_6443 : dirty_2_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7149 = _T_30 ? _GEN_6444 : dirty_2_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7150 = _T_30 ? _GEN_6445 : dirty_2_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7151 = _T_30 ? _GEN_6446 : dirty_2_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7152 = _T_30 ? _GEN_6447 : dirty_2_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7153 = _T_30 ? _GEN_6448 : dirty_2_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7154 = _T_30 ? _GEN_6449 : dirty_2_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7155 = _T_30 ? _GEN_6450 : dirty_2_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7156 = _T_30 ? _GEN_6451 : dirty_3_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7157 = _T_30 ? _GEN_6452 : dirty_3_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7158 = _T_30 ? _GEN_6453 : dirty_3_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7159 = _T_30 ? _GEN_6454 : dirty_3_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7160 = _T_30 ? _GEN_6455 : dirty_3_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7161 = _T_30 ? _GEN_6456 : dirty_3_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7162 = _T_30 ? _GEN_6457 : dirty_3_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7163 = _T_30 ? _GEN_6458 : dirty_3_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7164 = _T_30 ? _GEN_6459 : dirty_4_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7165 = _T_30 ? _GEN_6460 : dirty_4_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7166 = _T_30 ? _GEN_6461 : dirty_4_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7167 = _T_30 ? _GEN_6462 : dirty_4_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7168 = _T_30 ? _GEN_6463 : dirty_4_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7169 = _T_30 ? _GEN_6464 : dirty_4_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7170 = _T_30 ? _GEN_6465 : dirty_4_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7171 = _T_30 ? _GEN_6466 : dirty_4_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7172 = _T_30 ? _GEN_6467 : dirty_5_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7173 = _T_30 ? _GEN_6468 : dirty_5_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7174 = _T_30 ? _GEN_6469 : dirty_5_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7175 = _T_30 ? _GEN_6470 : dirty_5_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7176 = _T_30 ? _GEN_6471 : dirty_5_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7177 = _T_30 ? _GEN_6472 : dirty_5_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7178 = _T_30 ? _GEN_6473 : dirty_5_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7179 = _T_30 ? _GEN_6474 : dirty_5_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7180 = _T_30 ? _GEN_6475 : dirty_6_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7181 = _T_30 ? _GEN_6476 : dirty_6_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7182 = _T_30 ? _GEN_6477 : dirty_6_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7183 = _T_30 ? _GEN_6478 : dirty_6_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7184 = _T_30 ? _GEN_6479 : dirty_6_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7185 = _T_30 ? _GEN_6480 : dirty_6_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7186 = _T_30 ? _GEN_6481 : dirty_6_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7187 = _T_30 ? _GEN_6482 : dirty_6_7; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7188 = _T_30 ? _GEN_6483 : dirty_7_0; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7189 = _T_30 ? _GEN_6484 : dirty_7_1; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7190 = _T_30 ? _GEN_6485 : dirty_7_2; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7191 = _T_30 ? _GEN_6486 : dirty_7_3; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7192 = _T_30 ? _GEN_6487 : dirty_7_4; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7193 = _T_30 ? _GEN_6488 : dirty_7_5; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7194 = _T_30 ? _GEN_6489 : dirty_7_6; // @[Cache.scala 126:21 58:22]
  wire  _GEN_7195 = _T_30 ? _GEN_6490 : dirty_7_7; // @[Cache.scala 126:21 58:22]
  wire [31:0] _GEN_7196 = _T_30 ? _GEN_6491 : CacheMem_0_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7197 = _T_30 ? _GEN_6492 : CacheMem_0_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7198 = _T_30 ? _GEN_6493 : CacheMem_0_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7199 = _T_30 ? _GEN_6494 : CacheMem_0_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7200 = _T_30 ? _GEN_6495 : CacheMem_0_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7201 = _T_30 ? _GEN_6496 : CacheMem_0_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7202 = _T_30 ? _GEN_6497 : CacheMem_0_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7203 = _T_30 ? _GEN_6498 : CacheMem_0_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7204 = _T_30 ? _GEN_6499 : CacheMem_1_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7205 = _T_30 ? _GEN_6500 : CacheMem_1_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7206 = _T_30 ? _GEN_6501 : CacheMem_1_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7207 = _T_30 ? _GEN_6502 : CacheMem_1_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7208 = _T_30 ? _GEN_6503 : CacheMem_1_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7209 = _T_30 ? _GEN_6504 : CacheMem_1_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7210 = _T_30 ? _GEN_6505 : CacheMem_1_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7211 = _T_30 ? _GEN_6506 : CacheMem_1_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7212 = _T_30 ? _GEN_6507 : CacheMem_2_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7213 = _T_30 ? _GEN_6508 : CacheMem_2_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7214 = _T_30 ? _GEN_6509 : CacheMem_2_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7215 = _T_30 ? _GEN_6510 : CacheMem_2_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7216 = _T_30 ? _GEN_6511 : CacheMem_2_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7217 = _T_30 ? _GEN_6512 : CacheMem_2_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7218 = _T_30 ? _GEN_6513 : CacheMem_2_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7219 = _T_30 ? _GEN_6514 : CacheMem_2_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7220 = _T_30 ? _GEN_6515 : CacheMem_3_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7221 = _T_30 ? _GEN_6516 : CacheMem_3_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7222 = _T_30 ? _GEN_6517 : CacheMem_3_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7223 = _T_30 ? _GEN_6518 : CacheMem_3_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7224 = _T_30 ? _GEN_6519 : CacheMem_3_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7225 = _T_30 ? _GEN_6520 : CacheMem_3_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7226 = _T_30 ? _GEN_6521 : CacheMem_3_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7227 = _T_30 ? _GEN_6522 : CacheMem_3_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7228 = _T_30 ? _GEN_6523 : CacheMem_4_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7229 = _T_30 ? _GEN_6524 : CacheMem_4_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7230 = _T_30 ? _GEN_6525 : CacheMem_4_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7231 = _T_30 ? _GEN_6526 : CacheMem_4_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7232 = _T_30 ? _GEN_6527 : CacheMem_4_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7233 = _T_30 ? _GEN_6528 : CacheMem_4_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7234 = _T_30 ? _GEN_6529 : CacheMem_4_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7235 = _T_30 ? _GEN_6530 : CacheMem_4_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7236 = _T_30 ? _GEN_6531 : CacheMem_5_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7237 = _T_30 ? _GEN_6532 : CacheMem_5_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7238 = _T_30 ? _GEN_6533 : CacheMem_5_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7239 = _T_30 ? _GEN_6534 : CacheMem_5_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7240 = _T_30 ? _GEN_6535 : CacheMem_5_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7241 = _T_30 ? _GEN_6536 : CacheMem_5_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7242 = _T_30 ? _GEN_6537 : CacheMem_5_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7243 = _T_30 ? _GEN_6538 : CacheMem_5_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7244 = _T_30 ? _GEN_6539 : CacheMem_6_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7245 = _T_30 ? _GEN_6540 : CacheMem_6_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7246 = _T_30 ? _GEN_6541 : CacheMem_6_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7247 = _T_30 ? _GEN_6542 : CacheMem_6_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7248 = _T_30 ? _GEN_6543 : CacheMem_6_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7249 = _T_30 ? _GEN_6544 : CacheMem_6_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7250 = _T_30 ? _GEN_6545 : CacheMem_6_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7251 = _T_30 ? _GEN_6546 : CacheMem_6_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7252 = _T_30 ? _GEN_6547 : CacheMem_7_0_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7253 = _T_30 ? _GEN_6548 : CacheMem_7_1_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7254 = _T_30 ? _GEN_6549 : CacheMem_7_2_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7255 = _T_30 ? _GEN_6550 : CacheMem_7_3_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7256 = _T_30 ? _GEN_6551 : CacheMem_7_4_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7257 = _T_30 ? _GEN_6552 : CacheMem_7_5_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7258 = _T_30 ? _GEN_6553 : CacheMem_7_6_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7259 = _T_30 ? _GEN_6554 : CacheMem_7_7_0; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7260 = _T_30 ? _GEN_6555 : CacheMem_0_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7261 = _T_30 ? _GEN_6556 : CacheMem_0_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7262 = _T_30 ? _GEN_6557 : CacheMem_0_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7263 = _T_30 ? _GEN_6558 : CacheMem_0_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7264 = _T_30 ? _GEN_6559 : CacheMem_0_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7265 = _T_30 ? _GEN_6560 : CacheMem_0_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7266 = _T_30 ? _GEN_6561 : CacheMem_0_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7267 = _T_30 ? _GEN_6562 : CacheMem_0_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7268 = _T_30 ? _GEN_6563 : CacheMem_1_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7269 = _T_30 ? _GEN_6564 : CacheMem_1_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7270 = _T_30 ? _GEN_6565 : CacheMem_1_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7271 = _T_30 ? _GEN_6566 : CacheMem_1_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7272 = _T_30 ? _GEN_6567 : CacheMem_1_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7273 = _T_30 ? _GEN_6568 : CacheMem_1_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7274 = _T_30 ? _GEN_6569 : CacheMem_1_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7275 = _T_30 ? _GEN_6570 : CacheMem_1_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7276 = _T_30 ? _GEN_6571 : CacheMem_2_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7277 = _T_30 ? _GEN_6572 : CacheMem_2_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7278 = _T_30 ? _GEN_6573 : CacheMem_2_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7279 = _T_30 ? _GEN_6574 : CacheMem_2_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7280 = _T_30 ? _GEN_6575 : CacheMem_2_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7281 = _T_30 ? _GEN_6576 : CacheMem_2_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7282 = _T_30 ? _GEN_6577 : CacheMem_2_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7283 = _T_30 ? _GEN_6578 : CacheMem_2_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7284 = _T_30 ? _GEN_6579 : CacheMem_3_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7285 = _T_30 ? _GEN_6580 : CacheMem_3_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7286 = _T_30 ? _GEN_6581 : CacheMem_3_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7287 = _T_30 ? _GEN_6582 : CacheMem_3_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7288 = _T_30 ? _GEN_6583 : CacheMem_3_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7289 = _T_30 ? _GEN_6584 : CacheMem_3_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7290 = _T_30 ? _GEN_6585 : CacheMem_3_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7291 = _T_30 ? _GEN_6586 : CacheMem_3_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7292 = _T_30 ? _GEN_6587 : CacheMem_4_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7293 = _T_30 ? _GEN_6588 : CacheMem_4_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7294 = _T_30 ? _GEN_6589 : CacheMem_4_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7295 = _T_30 ? _GEN_6590 : CacheMem_4_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7296 = _T_30 ? _GEN_6591 : CacheMem_4_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7297 = _T_30 ? _GEN_6592 : CacheMem_4_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7298 = _T_30 ? _GEN_6593 : CacheMem_4_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7299 = _T_30 ? _GEN_6594 : CacheMem_4_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7300 = _T_30 ? _GEN_6595 : CacheMem_5_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7301 = _T_30 ? _GEN_6596 : CacheMem_5_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7302 = _T_30 ? _GEN_6597 : CacheMem_5_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7303 = _T_30 ? _GEN_6598 : CacheMem_5_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7304 = _T_30 ? _GEN_6599 : CacheMem_5_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7305 = _T_30 ? _GEN_6600 : CacheMem_5_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7306 = _T_30 ? _GEN_6601 : CacheMem_5_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7307 = _T_30 ? _GEN_6602 : CacheMem_5_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7308 = _T_30 ? _GEN_6603 : CacheMem_6_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7309 = _T_30 ? _GEN_6604 : CacheMem_6_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7310 = _T_30 ? _GEN_6605 : CacheMem_6_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7311 = _T_30 ? _GEN_6606 : CacheMem_6_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7312 = _T_30 ? _GEN_6607 : CacheMem_6_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7313 = _T_30 ? _GEN_6608 : CacheMem_6_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7314 = _T_30 ? _GEN_6609 : CacheMem_6_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7315 = _T_30 ? _GEN_6610 : CacheMem_6_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7316 = _T_30 ? _GEN_6611 : CacheMem_7_0_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7317 = _T_30 ? _GEN_6612 : CacheMem_7_1_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7318 = _T_30 ? _GEN_6613 : CacheMem_7_2_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7319 = _T_30 ? _GEN_6614 : CacheMem_7_3_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7320 = _T_30 ? _GEN_6615 : CacheMem_7_4_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7321 = _T_30 ? _GEN_6616 : CacheMem_7_5_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7322 = _T_30 ? _GEN_6617 : CacheMem_7_6_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7323 = _T_30 ? _GEN_6618 : CacheMem_7_7_1; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7324 = _T_30 ? _GEN_6619 : CacheMem_0_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7325 = _T_30 ? _GEN_6620 : CacheMem_0_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7326 = _T_30 ? _GEN_6621 : CacheMem_0_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7327 = _T_30 ? _GEN_6622 : CacheMem_0_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7328 = _T_30 ? _GEN_6623 : CacheMem_0_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7329 = _T_30 ? _GEN_6624 : CacheMem_0_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7330 = _T_30 ? _GEN_6625 : CacheMem_0_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7331 = _T_30 ? _GEN_6626 : CacheMem_0_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7332 = _T_30 ? _GEN_6627 : CacheMem_1_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7333 = _T_30 ? _GEN_6628 : CacheMem_1_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7334 = _T_30 ? _GEN_6629 : CacheMem_1_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7335 = _T_30 ? _GEN_6630 : CacheMem_1_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7336 = _T_30 ? _GEN_6631 : CacheMem_1_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7337 = _T_30 ? _GEN_6632 : CacheMem_1_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7338 = _T_30 ? _GEN_6633 : CacheMem_1_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7339 = _T_30 ? _GEN_6634 : CacheMem_1_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7340 = _T_30 ? _GEN_6635 : CacheMem_2_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7341 = _T_30 ? _GEN_6636 : CacheMem_2_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7342 = _T_30 ? _GEN_6637 : CacheMem_2_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7343 = _T_30 ? _GEN_6638 : CacheMem_2_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7344 = _T_30 ? _GEN_6639 : CacheMem_2_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7345 = _T_30 ? _GEN_6640 : CacheMem_2_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7346 = _T_30 ? _GEN_6641 : CacheMem_2_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7347 = _T_30 ? _GEN_6642 : CacheMem_2_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7348 = _T_30 ? _GEN_6643 : CacheMem_3_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7349 = _T_30 ? _GEN_6644 : CacheMem_3_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7350 = _T_30 ? _GEN_6645 : CacheMem_3_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7351 = _T_30 ? _GEN_6646 : CacheMem_3_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7352 = _T_30 ? _GEN_6647 : CacheMem_3_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7353 = _T_30 ? _GEN_6648 : CacheMem_3_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7354 = _T_30 ? _GEN_6649 : CacheMem_3_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7355 = _T_30 ? _GEN_6650 : CacheMem_3_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7356 = _T_30 ? _GEN_6651 : CacheMem_4_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7357 = _T_30 ? _GEN_6652 : CacheMem_4_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7358 = _T_30 ? _GEN_6653 : CacheMem_4_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7359 = _T_30 ? _GEN_6654 : CacheMem_4_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7360 = _T_30 ? _GEN_6655 : CacheMem_4_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7361 = _T_30 ? _GEN_6656 : CacheMem_4_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7362 = _T_30 ? _GEN_6657 : CacheMem_4_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7363 = _T_30 ? _GEN_6658 : CacheMem_4_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7364 = _T_30 ? _GEN_6659 : CacheMem_5_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7365 = _T_30 ? _GEN_6660 : CacheMem_5_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7366 = _T_30 ? _GEN_6661 : CacheMem_5_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7367 = _T_30 ? _GEN_6662 : CacheMem_5_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7368 = _T_30 ? _GEN_6663 : CacheMem_5_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7369 = _T_30 ? _GEN_6664 : CacheMem_5_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7370 = _T_30 ? _GEN_6665 : CacheMem_5_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7371 = _T_30 ? _GEN_6666 : CacheMem_5_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7372 = _T_30 ? _GEN_6667 : CacheMem_6_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7373 = _T_30 ? _GEN_6668 : CacheMem_6_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7374 = _T_30 ? _GEN_6669 : CacheMem_6_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7375 = _T_30 ? _GEN_6670 : CacheMem_6_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7376 = _T_30 ? _GEN_6671 : CacheMem_6_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7377 = _T_30 ? _GEN_6672 : CacheMem_6_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7378 = _T_30 ? _GEN_6673 : CacheMem_6_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7379 = _T_30 ? _GEN_6674 : CacheMem_6_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7380 = _T_30 ? _GEN_6675 : CacheMem_7_0_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7381 = _T_30 ? _GEN_6676 : CacheMem_7_1_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7382 = _T_30 ? _GEN_6677 : CacheMem_7_2_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7383 = _T_30 ? _GEN_6678 : CacheMem_7_3_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7384 = _T_30 ? _GEN_6679 : CacheMem_7_4_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7385 = _T_30 ? _GEN_6680 : CacheMem_7_5_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7386 = _T_30 ? _GEN_6681 : CacheMem_7_6_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7387 = _T_30 ? _GEN_6682 : CacheMem_7_7_2; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7388 = _T_30 ? _GEN_6683 : CacheMem_0_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7389 = _T_30 ? _GEN_6684 : CacheMem_0_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7390 = _T_30 ? _GEN_6685 : CacheMem_0_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7391 = _T_30 ? _GEN_6686 : CacheMem_0_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7392 = _T_30 ? _GEN_6687 : CacheMem_0_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7393 = _T_30 ? _GEN_6688 : CacheMem_0_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7394 = _T_30 ? _GEN_6689 : CacheMem_0_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7395 = _T_30 ? _GEN_6690 : CacheMem_0_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7396 = _T_30 ? _GEN_6691 : CacheMem_1_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7397 = _T_30 ? _GEN_6692 : CacheMem_1_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7398 = _T_30 ? _GEN_6693 : CacheMem_1_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7399 = _T_30 ? _GEN_6694 : CacheMem_1_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7400 = _T_30 ? _GEN_6695 : CacheMem_1_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7401 = _T_30 ? _GEN_6696 : CacheMem_1_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7402 = _T_30 ? _GEN_6697 : CacheMem_1_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7403 = _T_30 ? _GEN_6698 : CacheMem_1_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7404 = _T_30 ? _GEN_6699 : CacheMem_2_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7405 = _T_30 ? _GEN_6700 : CacheMem_2_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7406 = _T_30 ? _GEN_6701 : CacheMem_2_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7407 = _T_30 ? _GEN_6702 : CacheMem_2_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7408 = _T_30 ? _GEN_6703 : CacheMem_2_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7409 = _T_30 ? _GEN_6704 : CacheMem_2_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7410 = _T_30 ? _GEN_6705 : CacheMem_2_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7411 = _T_30 ? _GEN_6706 : CacheMem_2_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7412 = _T_30 ? _GEN_6707 : CacheMem_3_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7413 = _T_30 ? _GEN_6708 : CacheMem_3_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7414 = _T_30 ? _GEN_6709 : CacheMem_3_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7415 = _T_30 ? _GEN_6710 : CacheMem_3_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7416 = _T_30 ? _GEN_6711 : CacheMem_3_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7417 = _T_30 ? _GEN_6712 : CacheMem_3_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7418 = _T_30 ? _GEN_6713 : CacheMem_3_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7419 = _T_30 ? _GEN_6714 : CacheMem_3_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7420 = _T_30 ? _GEN_6715 : CacheMem_4_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7421 = _T_30 ? _GEN_6716 : CacheMem_4_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7422 = _T_30 ? _GEN_6717 : CacheMem_4_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7423 = _T_30 ? _GEN_6718 : CacheMem_4_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7424 = _T_30 ? _GEN_6719 : CacheMem_4_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7425 = _T_30 ? _GEN_6720 : CacheMem_4_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7426 = _T_30 ? _GEN_6721 : CacheMem_4_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7427 = _T_30 ? _GEN_6722 : CacheMem_4_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7428 = _T_30 ? _GEN_6723 : CacheMem_5_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7429 = _T_30 ? _GEN_6724 : CacheMem_5_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7430 = _T_30 ? _GEN_6725 : CacheMem_5_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7431 = _T_30 ? _GEN_6726 : CacheMem_5_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7432 = _T_30 ? _GEN_6727 : CacheMem_5_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7433 = _T_30 ? _GEN_6728 : CacheMem_5_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7434 = _T_30 ? _GEN_6729 : CacheMem_5_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7435 = _T_30 ? _GEN_6730 : CacheMem_5_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7436 = _T_30 ? _GEN_6731 : CacheMem_6_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7437 = _T_30 ? _GEN_6732 : CacheMem_6_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7438 = _T_30 ? _GEN_6733 : CacheMem_6_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7439 = _T_30 ? _GEN_6734 : CacheMem_6_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7440 = _T_30 ? _GEN_6735 : CacheMem_6_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7441 = _T_30 ? _GEN_6736 : CacheMem_6_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7442 = _T_30 ? _GEN_6737 : CacheMem_6_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7443 = _T_30 ? _GEN_6738 : CacheMem_6_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7444 = _T_30 ? _GEN_6739 : CacheMem_7_0_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7445 = _T_30 ? _GEN_6740 : CacheMem_7_1_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7446 = _T_30 ? _GEN_6741 : CacheMem_7_2_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7447 = _T_30 ? _GEN_6742 : CacheMem_7_3_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7448 = _T_30 ? _GEN_6743 : CacheMem_7_4_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7449 = _T_30 ? _GEN_6744 : CacheMem_7_5_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7450 = _T_30 ? _GEN_6745 : CacheMem_7_6_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7451 = _T_30 ? _GEN_6746 : CacheMem_7_7_3; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7452 = _T_30 ? _GEN_6747 : CacheMem_0_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7453 = _T_30 ? _GEN_6748 : CacheMem_0_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7454 = _T_30 ? _GEN_6749 : CacheMem_0_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7455 = _T_30 ? _GEN_6750 : CacheMem_0_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7456 = _T_30 ? _GEN_6751 : CacheMem_0_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7457 = _T_30 ? _GEN_6752 : CacheMem_0_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7458 = _T_30 ? _GEN_6753 : CacheMem_0_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7459 = _T_30 ? _GEN_6754 : CacheMem_0_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7460 = _T_30 ? _GEN_6755 : CacheMem_1_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7461 = _T_30 ? _GEN_6756 : CacheMem_1_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7462 = _T_30 ? _GEN_6757 : CacheMem_1_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7463 = _T_30 ? _GEN_6758 : CacheMem_1_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7464 = _T_30 ? _GEN_6759 : CacheMem_1_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7465 = _T_30 ? _GEN_6760 : CacheMem_1_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7466 = _T_30 ? _GEN_6761 : CacheMem_1_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7467 = _T_30 ? _GEN_6762 : CacheMem_1_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7468 = _T_30 ? _GEN_6763 : CacheMem_2_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7469 = _T_30 ? _GEN_6764 : CacheMem_2_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7470 = _T_30 ? _GEN_6765 : CacheMem_2_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7471 = _T_30 ? _GEN_6766 : CacheMem_2_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7472 = _T_30 ? _GEN_6767 : CacheMem_2_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7473 = _T_30 ? _GEN_6768 : CacheMem_2_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7474 = _T_30 ? _GEN_6769 : CacheMem_2_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7475 = _T_30 ? _GEN_6770 : CacheMem_2_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7476 = _T_30 ? _GEN_6771 : CacheMem_3_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7477 = _T_30 ? _GEN_6772 : CacheMem_3_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7478 = _T_30 ? _GEN_6773 : CacheMem_3_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7479 = _T_30 ? _GEN_6774 : CacheMem_3_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7480 = _T_30 ? _GEN_6775 : CacheMem_3_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7481 = _T_30 ? _GEN_6776 : CacheMem_3_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7482 = _T_30 ? _GEN_6777 : CacheMem_3_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7483 = _T_30 ? _GEN_6778 : CacheMem_3_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7484 = _T_30 ? _GEN_6779 : CacheMem_4_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7485 = _T_30 ? _GEN_6780 : CacheMem_4_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7486 = _T_30 ? _GEN_6781 : CacheMem_4_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7487 = _T_30 ? _GEN_6782 : CacheMem_4_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7488 = _T_30 ? _GEN_6783 : CacheMem_4_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7489 = _T_30 ? _GEN_6784 : CacheMem_4_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7490 = _T_30 ? _GEN_6785 : CacheMem_4_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7491 = _T_30 ? _GEN_6786 : CacheMem_4_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7492 = _T_30 ? _GEN_6787 : CacheMem_5_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7493 = _T_30 ? _GEN_6788 : CacheMem_5_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7494 = _T_30 ? _GEN_6789 : CacheMem_5_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7495 = _T_30 ? _GEN_6790 : CacheMem_5_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7496 = _T_30 ? _GEN_6791 : CacheMem_5_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7497 = _T_30 ? _GEN_6792 : CacheMem_5_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7498 = _T_30 ? _GEN_6793 : CacheMem_5_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7499 = _T_30 ? _GEN_6794 : CacheMem_5_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7500 = _T_30 ? _GEN_6795 : CacheMem_6_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7501 = _T_30 ? _GEN_6796 : CacheMem_6_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7502 = _T_30 ? _GEN_6797 : CacheMem_6_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7503 = _T_30 ? _GEN_6798 : CacheMem_6_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7504 = _T_30 ? _GEN_6799 : CacheMem_6_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7505 = _T_30 ? _GEN_6800 : CacheMem_6_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7506 = _T_30 ? _GEN_6801 : CacheMem_6_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7507 = _T_30 ? _GEN_6802 : CacheMem_6_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7508 = _T_30 ? _GEN_6803 : CacheMem_7_0_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7509 = _T_30 ? _GEN_6804 : CacheMem_7_1_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7510 = _T_30 ? _GEN_6805 : CacheMem_7_2_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7511 = _T_30 ? _GEN_6806 : CacheMem_7_3_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7512 = _T_30 ? _GEN_6807 : CacheMem_7_4_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7513 = _T_30 ? _GEN_6808 : CacheMem_7_5_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7514 = _T_30 ? _GEN_6809 : CacheMem_7_6_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7515 = _T_30 ? _GEN_6810 : CacheMem_7_7_4; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7516 = _T_30 ? _GEN_6811 : CacheMem_0_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7517 = _T_30 ? _GEN_6812 : CacheMem_0_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7518 = _T_30 ? _GEN_6813 : CacheMem_0_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7519 = _T_30 ? _GEN_6814 : CacheMem_0_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7520 = _T_30 ? _GEN_6815 : CacheMem_0_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7521 = _T_30 ? _GEN_6816 : CacheMem_0_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7522 = _T_30 ? _GEN_6817 : CacheMem_0_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7523 = _T_30 ? _GEN_6818 : CacheMem_0_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7524 = _T_30 ? _GEN_6819 : CacheMem_1_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7525 = _T_30 ? _GEN_6820 : CacheMem_1_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7526 = _T_30 ? _GEN_6821 : CacheMem_1_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7527 = _T_30 ? _GEN_6822 : CacheMem_1_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7528 = _T_30 ? _GEN_6823 : CacheMem_1_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7529 = _T_30 ? _GEN_6824 : CacheMem_1_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7530 = _T_30 ? _GEN_6825 : CacheMem_1_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7531 = _T_30 ? _GEN_6826 : CacheMem_1_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7532 = _T_30 ? _GEN_6827 : CacheMem_2_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7533 = _T_30 ? _GEN_6828 : CacheMem_2_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7534 = _T_30 ? _GEN_6829 : CacheMem_2_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7535 = _T_30 ? _GEN_6830 : CacheMem_2_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7536 = _T_30 ? _GEN_6831 : CacheMem_2_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7537 = _T_30 ? _GEN_6832 : CacheMem_2_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7538 = _T_30 ? _GEN_6833 : CacheMem_2_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7539 = _T_30 ? _GEN_6834 : CacheMem_2_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7540 = _T_30 ? _GEN_6835 : CacheMem_3_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7541 = _T_30 ? _GEN_6836 : CacheMem_3_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7542 = _T_30 ? _GEN_6837 : CacheMem_3_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7543 = _T_30 ? _GEN_6838 : CacheMem_3_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7544 = _T_30 ? _GEN_6839 : CacheMem_3_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7545 = _T_30 ? _GEN_6840 : CacheMem_3_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7546 = _T_30 ? _GEN_6841 : CacheMem_3_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7547 = _T_30 ? _GEN_6842 : CacheMem_3_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7548 = _T_30 ? _GEN_6843 : CacheMem_4_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7549 = _T_30 ? _GEN_6844 : CacheMem_4_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7550 = _T_30 ? _GEN_6845 : CacheMem_4_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7551 = _T_30 ? _GEN_6846 : CacheMem_4_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7552 = _T_30 ? _GEN_6847 : CacheMem_4_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7553 = _T_30 ? _GEN_6848 : CacheMem_4_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7554 = _T_30 ? _GEN_6849 : CacheMem_4_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7555 = _T_30 ? _GEN_6850 : CacheMem_4_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7556 = _T_30 ? _GEN_6851 : CacheMem_5_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7557 = _T_30 ? _GEN_6852 : CacheMem_5_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7558 = _T_30 ? _GEN_6853 : CacheMem_5_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7559 = _T_30 ? _GEN_6854 : CacheMem_5_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7560 = _T_30 ? _GEN_6855 : CacheMem_5_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7561 = _T_30 ? _GEN_6856 : CacheMem_5_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7562 = _T_30 ? _GEN_6857 : CacheMem_5_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7563 = _T_30 ? _GEN_6858 : CacheMem_5_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7564 = _T_30 ? _GEN_6859 : CacheMem_6_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7565 = _T_30 ? _GEN_6860 : CacheMem_6_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7566 = _T_30 ? _GEN_6861 : CacheMem_6_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7567 = _T_30 ? _GEN_6862 : CacheMem_6_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7568 = _T_30 ? _GEN_6863 : CacheMem_6_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7569 = _T_30 ? _GEN_6864 : CacheMem_6_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7570 = _T_30 ? _GEN_6865 : CacheMem_6_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7571 = _T_30 ? _GEN_6866 : CacheMem_6_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7572 = _T_30 ? _GEN_6867 : CacheMem_7_0_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7573 = _T_30 ? _GEN_6868 : CacheMem_7_1_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7574 = _T_30 ? _GEN_6869 : CacheMem_7_2_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7575 = _T_30 ? _GEN_6870 : CacheMem_7_3_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7576 = _T_30 ? _GEN_6871 : CacheMem_7_4_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7577 = _T_30 ? _GEN_6872 : CacheMem_7_5_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7578 = _T_30 ? _GEN_6873 : CacheMem_7_6_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7579 = _T_30 ? _GEN_6874 : CacheMem_7_7_5; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7580 = _T_30 ? _GEN_6875 : CacheMem_0_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7581 = _T_30 ? _GEN_6876 : CacheMem_0_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7582 = _T_30 ? _GEN_6877 : CacheMem_0_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7583 = _T_30 ? _GEN_6878 : CacheMem_0_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7584 = _T_30 ? _GEN_6879 : CacheMem_0_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7585 = _T_30 ? _GEN_6880 : CacheMem_0_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7586 = _T_30 ? _GEN_6881 : CacheMem_0_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7587 = _T_30 ? _GEN_6882 : CacheMem_0_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7588 = _T_30 ? _GEN_6883 : CacheMem_1_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7589 = _T_30 ? _GEN_6884 : CacheMem_1_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7590 = _T_30 ? _GEN_6885 : CacheMem_1_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7591 = _T_30 ? _GEN_6886 : CacheMem_1_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7592 = _T_30 ? _GEN_6887 : CacheMem_1_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7593 = _T_30 ? _GEN_6888 : CacheMem_1_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7594 = _T_30 ? _GEN_6889 : CacheMem_1_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7595 = _T_30 ? _GEN_6890 : CacheMem_1_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7596 = _T_30 ? _GEN_6891 : CacheMem_2_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7597 = _T_30 ? _GEN_6892 : CacheMem_2_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7598 = _T_30 ? _GEN_6893 : CacheMem_2_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7599 = _T_30 ? _GEN_6894 : CacheMem_2_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7600 = _T_30 ? _GEN_6895 : CacheMem_2_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7601 = _T_30 ? _GEN_6896 : CacheMem_2_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7602 = _T_30 ? _GEN_6897 : CacheMem_2_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7603 = _T_30 ? _GEN_6898 : CacheMem_2_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7604 = _T_30 ? _GEN_6899 : CacheMem_3_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7605 = _T_30 ? _GEN_6900 : CacheMem_3_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7606 = _T_30 ? _GEN_6901 : CacheMem_3_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7607 = _T_30 ? _GEN_6902 : CacheMem_3_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7608 = _T_30 ? _GEN_6903 : CacheMem_3_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7609 = _T_30 ? _GEN_6904 : CacheMem_3_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7610 = _T_30 ? _GEN_6905 : CacheMem_3_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7611 = _T_30 ? _GEN_6906 : CacheMem_3_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7612 = _T_30 ? _GEN_6907 : CacheMem_4_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7613 = _T_30 ? _GEN_6908 : CacheMem_4_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7614 = _T_30 ? _GEN_6909 : CacheMem_4_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7615 = _T_30 ? _GEN_6910 : CacheMem_4_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7616 = _T_30 ? _GEN_6911 : CacheMem_4_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7617 = _T_30 ? _GEN_6912 : CacheMem_4_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7618 = _T_30 ? _GEN_6913 : CacheMem_4_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7619 = _T_30 ? _GEN_6914 : CacheMem_4_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7620 = _T_30 ? _GEN_6915 : CacheMem_5_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7621 = _T_30 ? _GEN_6916 : CacheMem_5_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7622 = _T_30 ? _GEN_6917 : CacheMem_5_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7623 = _T_30 ? _GEN_6918 : CacheMem_5_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7624 = _T_30 ? _GEN_6919 : CacheMem_5_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7625 = _T_30 ? _GEN_6920 : CacheMem_5_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7626 = _T_30 ? _GEN_6921 : CacheMem_5_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7627 = _T_30 ? _GEN_6922 : CacheMem_5_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7628 = _T_30 ? _GEN_6923 : CacheMem_6_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7629 = _T_30 ? _GEN_6924 : CacheMem_6_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7630 = _T_30 ? _GEN_6925 : CacheMem_6_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7631 = _T_30 ? _GEN_6926 : CacheMem_6_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7632 = _T_30 ? _GEN_6927 : CacheMem_6_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7633 = _T_30 ? _GEN_6928 : CacheMem_6_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7634 = _T_30 ? _GEN_6929 : CacheMem_6_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7635 = _T_30 ? _GEN_6930 : CacheMem_6_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7636 = _T_30 ? _GEN_6931 : CacheMem_7_0_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7637 = _T_30 ? _GEN_6932 : CacheMem_7_1_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7638 = _T_30 ? _GEN_6933 : CacheMem_7_2_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7639 = _T_30 ? _GEN_6934 : CacheMem_7_3_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7640 = _T_30 ? _GEN_6935 : CacheMem_7_4_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7641 = _T_30 ? _GEN_6936 : CacheMem_7_5_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7642 = _T_30 ? _GEN_6937 : CacheMem_7_6_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7643 = _T_30 ? _GEN_6938 : CacheMem_7_7_6; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7644 = _T_30 ? _GEN_6939 : CacheMem_0_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7645 = _T_30 ? _GEN_6940 : CacheMem_0_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7646 = _T_30 ? _GEN_6941 : CacheMem_0_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7647 = _T_30 ? _GEN_6942 : CacheMem_0_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7648 = _T_30 ? _GEN_6943 : CacheMem_0_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7649 = _T_30 ? _GEN_6944 : CacheMem_0_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7650 = _T_30 ? _GEN_6945 : CacheMem_0_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7651 = _T_30 ? _GEN_6946 : CacheMem_0_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7652 = _T_30 ? _GEN_6947 : CacheMem_1_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7653 = _T_30 ? _GEN_6948 : CacheMem_1_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7654 = _T_30 ? _GEN_6949 : CacheMem_1_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7655 = _T_30 ? _GEN_6950 : CacheMem_1_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7656 = _T_30 ? _GEN_6951 : CacheMem_1_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7657 = _T_30 ? _GEN_6952 : CacheMem_1_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7658 = _T_30 ? _GEN_6953 : CacheMem_1_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7659 = _T_30 ? _GEN_6954 : CacheMem_1_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7660 = _T_30 ? _GEN_6955 : CacheMem_2_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7661 = _T_30 ? _GEN_6956 : CacheMem_2_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7662 = _T_30 ? _GEN_6957 : CacheMem_2_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7663 = _T_30 ? _GEN_6958 : CacheMem_2_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7664 = _T_30 ? _GEN_6959 : CacheMem_2_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7665 = _T_30 ? _GEN_6960 : CacheMem_2_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7666 = _T_30 ? _GEN_6961 : CacheMem_2_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7667 = _T_30 ? _GEN_6962 : CacheMem_2_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7668 = _T_30 ? _GEN_6963 : CacheMem_3_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7669 = _T_30 ? _GEN_6964 : CacheMem_3_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7670 = _T_30 ? _GEN_6965 : CacheMem_3_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7671 = _T_30 ? _GEN_6966 : CacheMem_3_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7672 = _T_30 ? _GEN_6967 : CacheMem_3_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7673 = _T_30 ? _GEN_6968 : CacheMem_3_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7674 = _T_30 ? _GEN_6969 : CacheMem_3_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7675 = _T_30 ? _GEN_6970 : CacheMem_3_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7676 = _T_30 ? _GEN_6971 : CacheMem_4_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7677 = _T_30 ? _GEN_6972 : CacheMem_4_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7678 = _T_30 ? _GEN_6973 : CacheMem_4_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7679 = _T_30 ? _GEN_6974 : CacheMem_4_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7680 = _T_30 ? _GEN_6975 : CacheMem_4_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7681 = _T_30 ? _GEN_6976 : CacheMem_4_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7682 = _T_30 ? _GEN_6977 : CacheMem_4_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7683 = _T_30 ? _GEN_6978 : CacheMem_4_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7684 = _T_30 ? _GEN_6979 : CacheMem_5_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7685 = _T_30 ? _GEN_6980 : CacheMem_5_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7686 = _T_30 ? _GEN_6981 : CacheMem_5_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7687 = _T_30 ? _GEN_6982 : CacheMem_5_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7688 = _T_30 ? _GEN_6983 : CacheMem_5_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7689 = _T_30 ? _GEN_6984 : CacheMem_5_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7690 = _T_30 ? _GEN_6985 : CacheMem_5_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7691 = _T_30 ? _GEN_6986 : CacheMem_5_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7692 = _T_30 ? _GEN_6987 : CacheMem_6_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7693 = _T_30 ? _GEN_6988 : CacheMem_6_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7694 = _T_30 ? _GEN_6989 : CacheMem_6_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7695 = _T_30 ? _GEN_6990 : CacheMem_6_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7696 = _T_30 ? _GEN_6991 : CacheMem_6_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7697 = _T_30 ? _GEN_6992 : CacheMem_6_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7698 = _T_30 ? _GEN_6993 : CacheMem_6_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7699 = _T_30 ? _GEN_6994 : CacheMem_6_7_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7700 = _T_30 ? _GEN_6995 : CacheMem_7_0_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7701 = _T_30 ? _GEN_6996 : CacheMem_7_1_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7702 = _T_30 ? _GEN_6997 : CacheMem_7_2_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7703 = _T_30 ? _GEN_6998 : CacheMem_7_3_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7704 = _T_30 ? _GEN_6999 : CacheMem_7_4_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7705 = _T_30 ? _GEN_7000 : CacheMem_7_5_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7706 = _T_30 ? _GEN_7001 : CacheMem_7_6_7; // @[Cache.scala 126:21 53:25]
  wire [31:0] _GEN_7707 = _T_30 ? _GEN_7002 : CacheMem_7_7_7; // @[Cache.scala 126:21 53:25]
  wire [8:0] _io_mem_addr_T_1 = io_mem_wr_req ? mem_wr_addr : 9'h0; // @[Cache.scala 191:64]
  assign io_outdata = _T_27 ? _GEN_5708 : 32'h0; // @[Cache.scala 126:21]
  assign io_miss = (io_r_req | io_w_req) & ~(cache_Hit & cacheState == 2'h0); // @[Cache.scala 196:36]
  assign io_mem_addr = io_mem_rd_req ? mem_rd_addr : _io_mem_addr_T_1; // @[Cache.scala 191:21]
  assign io_mem_rd_req = cacheState == 2'h2; // @[Cache.scala 187:35]
  assign io_mem_wr_req = cacheState == 2'h1; // @[Cache.scala 188:35]
  assign io_mem_wr_line_0 = mem_wr_line_0; // @[Cache.scala 195:18]
  assign io_mem_wr_line_1 = mem_wr_line_1; // @[Cache.scala 195:18]
  assign io_mem_wr_line_2 = mem_wr_line_2; // @[Cache.scala 195:18]
  assign io_mem_wr_line_3 = mem_wr_line_3; // @[Cache.scala 195:18]
  assign io_mem_wr_line_4 = mem_wr_line_4; // @[Cache.scala 195:18]
  assign io_mem_wr_line_5 = mem_wr_line_5; // @[Cache.scala 195:18]
  assign io_mem_wr_line_6 = mem_wr_line_6; // @[Cache.scala 195:18]
  assign io_mem_wr_line_7 = mem_wr_line_7; // @[Cache.scala 195:18]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_0 <= _GEN_3827;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_0 <= _GEN_7196;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_1 <= _GEN_3828;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_1 <= _GEN_7260;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_2 <= _GEN_3829;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_2 <= _GEN_7324;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_3 <= _GEN_3830;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_3 <= _GEN_7388;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_4 <= _GEN_3831;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_4 <= _GEN_7452;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_5 <= _GEN_3832;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_5 <= _GEN_7516;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_6 <= _GEN_3833;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_6 <= _GEN_7580;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_0_7 <= _GEN_3834;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_0_7 <= _GEN_7644;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_0 <= _GEN_3835;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_0 <= _GEN_7197;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_1 <= _GEN_3836;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_1 <= _GEN_7261;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_2 <= _GEN_3837;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_2 <= _GEN_7325;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_3 <= _GEN_3838;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_3 <= _GEN_7389;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_4 <= _GEN_3839;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_4 <= _GEN_7453;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_5 <= _GEN_3840;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_5 <= _GEN_7517;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_6 <= _GEN_3841;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_6 <= _GEN_7581;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_1_7 <= _GEN_3842;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_1_7 <= _GEN_7645;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_0 <= _GEN_3843;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_0 <= _GEN_7198;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_1 <= _GEN_3844;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_1 <= _GEN_7262;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_2 <= _GEN_3845;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_2 <= _GEN_7326;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_3 <= _GEN_3846;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_3 <= _GEN_7390;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_4 <= _GEN_3847;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_4 <= _GEN_7454;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_5 <= _GEN_3848;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_5 <= _GEN_7518;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_6 <= _GEN_3849;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_6 <= _GEN_7582;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_2_7 <= _GEN_3850;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_2_7 <= _GEN_7646;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_0 <= _GEN_3851;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_0 <= _GEN_7199;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_1 <= _GEN_3852;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_1 <= _GEN_7263;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_2 <= _GEN_3853;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_2 <= _GEN_7327;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_3 <= _GEN_3854;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_3 <= _GEN_7391;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_4 <= _GEN_3855;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_4 <= _GEN_7455;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_5 <= _GEN_3856;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_5 <= _GEN_7519;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_6 <= _GEN_3857;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_6 <= _GEN_7583;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_3_7 <= _GEN_3858;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_3_7 <= _GEN_7647;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_0 <= _GEN_3859;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_0 <= _GEN_7200;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_1 <= _GEN_3860;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_1 <= _GEN_7264;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_2 <= _GEN_3861;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_2 <= _GEN_7328;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_3 <= _GEN_3862;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_3 <= _GEN_7392;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_4 <= _GEN_3863;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_4 <= _GEN_7456;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_5 <= _GEN_3864;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_5 <= _GEN_7520;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_6 <= _GEN_3865;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_6 <= _GEN_7584;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_4_7 <= _GEN_3866;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_4_7 <= _GEN_7648;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_0 <= _GEN_3867;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_0 <= _GEN_7201;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_1 <= _GEN_3868;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_1 <= _GEN_7265;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_2 <= _GEN_3869;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_2 <= _GEN_7329;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_3 <= _GEN_3870;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_3 <= _GEN_7393;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_4 <= _GEN_3871;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_4 <= _GEN_7457;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_5 <= _GEN_3872;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_5 <= _GEN_7521;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_6 <= _GEN_3873;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_6 <= _GEN_7585;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_5_7 <= _GEN_3874;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_5_7 <= _GEN_7649;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_0 <= _GEN_3875;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_0 <= _GEN_7202;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_1 <= _GEN_3876;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_1 <= _GEN_7266;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_2 <= _GEN_3877;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_2 <= _GEN_7330;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_3 <= _GEN_3878;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_3 <= _GEN_7394;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_4 <= _GEN_3879;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_4 <= _GEN_7458;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_5 <= _GEN_3880;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_5 <= _GEN_7522;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_6 <= _GEN_3881;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_6 <= _GEN_7586;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_6_7 <= _GEN_3882;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_6_7 <= _GEN_7650;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_0 <= _GEN_3883;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_0 <= _GEN_7203;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_1 <= _GEN_3884;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_1 <= _GEN_7267;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_2 <= _GEN_3885;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_2 <= _GEN_7331;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_3 <= _GEN_3886;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_3 <= _GEN_7395;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_4 <= _GEN_3887;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_4 <= _GEN_7459;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_5 <= _GEN_3888;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_5 <= _GEN_7523;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_6 <= _GEN_3889;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_6 <= _GEN_7587;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_0_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_0_7_7 <= _GEN_3890;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_0_7_7 <= _GEN_7651;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_0 <= _GEN_3891;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_0 <= _GEN_7204;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_1 <= _GEN_3892;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_1 <= _GEN_7268;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_2 <= _GEN_3893;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_2 <= _GEN_7332;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_3 <= _GEN_3894;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_3 <= _GEN_7396;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_4 <= _GEN_3895;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_4 <= _GEN_7460;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_5 <= _GEN_3896;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_5 <= _GEN_7524;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_6 <= _GEN_3897;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_6 <= _GEN_7588;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_0_7 <= _GEN_3898;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_0_7 <= _GEN_7652;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_0 <= _GEN_3899;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_0 <= _GEN_7205;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_1 <= _GEN_3900;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_1 <= _GEN_7269;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_2 <= _GEN_3901;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_2 <= _GEN_7333;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_3 <= _GEN_3902;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_3 <= _GEN_7397;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_4 <= _GEN_3903;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_4 <= _GEN_7461;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_5 <= _GEN_3904;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_5 <= _GEN_7525;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_6 <= _GEN_3905;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_6 <= _GEN_7589;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_1_7 <= _GEN_3906;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_1_7 <= _GEN_7653;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_0 <= _GEN_3907;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_0 <= _GEN_7206;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_1 <= _GEN_3908;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_1 <= _GEN_7270;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_2 <= _GEN_3909;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_2 <= _GEN_7334;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_3 <= _GEN_3910;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_3 <= _GEN_7398;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_4 <= _GEN_3911;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_4 <= _GEN_7462;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_5 <= _GEN_3912;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_5 <= _GEN_7526;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_6 <= _GEN_3913;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_6 <= _GEN_7590;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_2_7 <= _GEN_3914;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_2_7 <= _GEN_7654;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_0 <= _GEN_3915;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_0 <= _GEN_7207;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_1 <= _GEN_3916;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_1 <= _GEN_7271;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_2 <= _GEN_3917;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_2 <= _GEN_7335;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_3 <= _GEN_3918;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_3 <= _GEN_7399;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_4 <= _GEN_3919;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_4 <= _GEN_7463;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_5 <= _GEN_3920;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_5 <= _GEN_7527;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_6 <= _GEN_3921;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_6 <= _GEN_7591;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_3_7 <= _GEN_3922;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_3_7 <= _GEN_7655;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_0 <= _GEN_3923;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_0 <= _GEN_7208;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_1 <= _GEN_3924;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_1 <= _GEN_7272;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_2 <= _GEN_3925;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_2 <= _GEN_7336;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_3 <= _GEN_3926;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_3 <= _GEN_7400;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_4 <= _GEN_3927;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_4 <= _GEN_7464;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_5 <= _GEN_3928;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_5 <= _GEN_7528;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_6 <= _GEN_3929;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_6 <= _GEN_7592;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_4_7 <= _GEN_3930;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_4_7 <= _GEN_7656;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_0 <= _GEN_3931;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_0 <= _GEN_7209;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_1 <= _GEN_3932;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_1 <= _GEN_7273;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_2 <= _GEN_3933;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_2 <= _GEN_7337;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_3 <= _GEN_3934;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_3 <= _GEN_7401;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_4 <= _GEN_3935;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_4 <= _GEN_7465;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_5 <= _GEN_3936;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_5 <= _GEN_7529;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_6 <= _GEN_3937;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_6 <= _GEN_7593;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_5_7 <= _GEN_3938;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_5_7 <= _GEN_7657;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_0 <= _GEN_3939;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_0 <= _GEN_7210;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_1 <= _GEN_3940;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_1 <= _GEN_7274;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_2 <= _GEN_3941;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_2 <= _GEN_7338;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_3 <= _GEN_3942;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_3 <= _GEN_7402;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_4 <= _GEN_3943;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_4 <= _GEN_7466;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_5 <= _GEN_3944;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_5 <= _GEN_7530;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_6 <= _GEN_3945;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_6 <= _GEN_7594;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_6_7 <= _GEN_3946;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_6_7 <= _GEN_7658;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_0 <= _GEN_3947;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_0 <= _GEN_7211;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_1 <= _GEN_3948;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_1 <= _GEN_7275;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_2 <= _GEN_3949;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_2 <= _GEN_7339;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_3 <= _GEN_3950;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_3 <= _GEN_7403;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_4 <= _GEN_3951;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_4 <= _GEN_7467;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_5 <= _GEN_3952;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_5 <= _GEN_7531;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_6 <= _GEN_3953;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_6 <= _GEN_7595;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_1_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_1_7_7 <= _GEN_3954;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_1_7_7 <= _GEN_7659;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_0 <= _GEN_3955;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_0 <= _GEN_7212;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_1 <= _GEN_3956;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_1 <= _GEN_7276;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_2 <= _GEN_3957;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_2 <= _GEN_7340;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_3 <= _GEN_3958;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_3 <= _GEN_7404;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_4 <= _GEN_3959;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_4 <= _GEN_7468;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_5 <= _GEN_3960;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_5 <= _GEN_7532;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_6 <= _GEN_3961;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_6 <= _GEN_7596;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_0_7 <= _GEN_3962;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_0_7 <= _GEN_7660;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_0 <= _GEN_3963;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_0 <= _GEN_7213;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_1 <= _GEN_3964;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_1 <= _GEN_7277;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_2 <= _GEN_3965;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_2 <= _GEN_7341;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_3 <= _GEN_3966;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_3 <= _GEN_7405;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_4 <= _GEN_3967;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_4 <= _GEN_7469;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_5 <= _GEN_3968;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_5 <= _GEN_7533;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_6 <= _GEN_3969;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_6 <= _GEN_7597;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_1_7 <= _GEN_3970;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_1_7 <= _GEN_7661;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_0 <= _GEN_3971;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_0 <= _GEN_7214;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_1 <= _GEN_3972;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_1 <= _GEN_7278;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_2 <= _GEN_3973;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_2 <= _GEN_7342;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_3 <= _GEN_3974;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_3 <= _GEN_7406;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_4 <= _GEN_3975;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_4 <= _GEN_7470;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_5 <= _GEN_3976;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_5 <= _GEN_7534;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_6 <= _GEN_3977;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_6 <= _GEN_7598;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_2_7 <= _GEN_3978;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_2_7 <= _GEN_7662;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_0 <= _GEN_3979;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_0 <= _GEN_7215;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_1 <= _GEN_3980;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_1 <= _GEN_7279;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_2 <= _GEN_3981;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_2 <= _GEN_7343;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_3 <= _GEN_3982;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_3 <= _GEN_7407;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_4 <= _GEN_3983;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_4 <= _GEN_7471;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_5 <= _GEN_3984;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_5 <= _GEN_7535;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_6 <= _GEN_3985;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_6 <= _GEN_7599;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_3_7 <= _GEN_3986;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_3_7 <= _GEN_7663;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_0 <= _GEN_3987;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_0 <= _GEN_7216;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_1 <= _GEN_3988;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_1 <= _GEN_7280;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_2 <= _GEN_3989;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_2 <= _GEN_7344;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_3 <= _GEN_3990;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_3 <= _GEN_7408;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_4 <= _GEN_3991;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_4 <= _GEN_7472;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_5 <= _GEN_3992;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_5 <= _GEN_7536;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_6 <= _GEN_3993;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_6 <= _GEN_7600;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_4_7 <= _GEN_3994;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_4_7 <= _GEN_7664;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_0 <= _GEN_3995;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_0 <= _GEN_7217;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_1 <= _GEN_3996;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_1 <= _GEN_7281;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_2 <= _GEN_3997;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_2 <= _GEN_7345;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_3 <= _GEN_3998;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_3 <= _GEN_7409;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_4 <= _GEN_3999;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_4 <= _GEN_7473;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_5 <= _GEN_4000;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_5 <= _GEN_7537;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_6 <= _GEN_4001;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_6 <= _GEN_7601;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_5_7 <= _GEN_4002;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_5_7 <= _GEN_7665;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_0 <= _GEN_4003;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_0 <= _GEN_7218;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_1 <= _GEN_4004;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_1 <= _GEN_7282;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_2 <= _GEN_4005;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_2 <= _GEN_7346;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_3 <= _GEN_4006;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_3 <= _GEN_7410;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_4 <= _GEN_4007;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_4 <= _GEN_7474;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_5 <= _GEN_4008;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_5 <= _GEN_7538;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_6 <= _GEN_4009;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_6 <= _GEN_7602;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_6_7 <= _GEN_4010;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_6_7 <= _GEN_7666;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_0 <= _GEN_4011;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_0 <= _GEN_7219;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_1 <= _GEN_4012;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_1 <= _GEN_7283;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_2 <= _GEN_4013;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_2 <= _GEN_7347;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_3 <= _GEN_4014;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_3 <= _GEN_7411;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_4 <= _GEN_4015;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_4 <= _GEN_7475;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_5 <= _GEN_4016;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_5 <= _GEN_7539;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_6 <= _GEN_4017;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_6 <= _GEN_7603;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_2_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_2_7_7 <= _GEN_4018;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_2_7_7 <= _GEN_7667;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_0 <= _GEN_4019;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_0 <= _GEN_7220;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_1 <= _GEN_4020;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_1 <= _GEN_7284;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_2 <= _GEN_4021;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_2 <= _GEN_7348;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_3 <= _GEN_4022;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_3 <= _GEN_7412;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_4 <= _GEN_4023;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_4 <= _GEN_7476;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_5 <= _GEN_4024;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_5 <= _GEN_7540;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_6 <= _GEN_4025;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_6 <= _GEN_7604;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_0_7 <= _GEN_4026;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_0_7 <= _GEN_7668;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_0 <= _GEN_4027;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_0 <= _GEN_7221;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_1 <= _GEN_4028;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_1 <= _GEN_7285;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_2 <= _GEN_4029;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_2 <= _GEN_7349;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_3 <= _GEN_4030;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_3 <= _GEN_7413;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_4 <= _GEN_4031;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_4 <= _GEN_7477;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_5 <= _GEN_4032;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_5 <= _GEN_7541;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_6 <= _GEN_4033;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_6 <= _GEN_7605;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_1_7 <= _GEN_4034;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_1_7 <= _GEN_7669;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_0 <= _GEN_4035;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_0 <= _GEN_7222;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_1 <= _GEN_4036;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_1 <= _GEN_7286;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_2 <= _GEN_4037;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_2 <= _GEN_7350;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_3 <= _GEN_4038;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_3 <= _GEN_7414;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_4 <= _GEN_4039;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_4 <= _GEN_7478;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_5 <= _GEN_4040;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_5 <= _GEN_7542;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_6 <= _GEN_4041;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_6 <= _GEN_7606;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_2_7 <= _GEN_4042;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_2_7 <= _GEN_7670;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_0 <= _GEN_4043;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_0 <= _GEN_7223;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_1 <= _GEN_4044;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_1 <= _GEN_7287;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_2 <= _GEN_4045;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_2 <= _GEN_7351;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_3 <= _GEN_4046;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_3 <= _GEN_7415;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_4 <= _GEN_4047;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_4 <= _GEN_7479;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_5 <= _GEN_4048;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_5 <= _GEN_7543;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_6 <= _GEN_4049;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_6 <= _GEN_7607;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_3_7 <= _GEN_4050;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_3_7 <= _GEN_7671;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_0 <= _GEN_4051;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_0 <= _GEN_7224;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_1 <= _GEN_4052;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_1 <= _GEN_7288;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_2 <= _GEN_4053;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_2 <= _GEN_7352;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_3 <= _GEN_4054;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_3 <= _GEN_7416;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_4 <= _GEN_4055;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_4 <= _GEN_7480;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_5 <= _GEN_4056;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_5 <= _GEN_7544;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_6 <= _GEN_4057;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_6 <= _GEN_7608;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_4_7 <= _GEN_4058;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_4_7 <= _GEN_7672;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_0 <= _GEN_4059;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_0 <= _GEN_7225;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_1 <= _GEN_4060;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_1 <= _GEN_7289;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_2 <= _GEN_4061;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_2 <= _GEN_7353;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_3 <= _GEN_4062;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_3 <= _GEN_7417;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_4 <= _GEN_4063;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_4 <= _GEN_7481;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_5 <= _GEN_4064;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_5 <= _GEN_7545;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_6 <= _GEN_4065;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_6 <= _GEN_7609;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_5_7 <= _GEN_4066;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_5_7 <= _GEN_7673;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_0 <= _GEN_4067;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_0 <= _GEN_7226;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_1 <= _GEN_4068;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_1 <= _GEN_7290;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_2 <= _GEN_4069;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_2 <= _GEN_7354;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_3 <= _GEN_4070;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_3 <= _GEN_7418;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_4 <= _GEN_4071;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_4 <= _GEN_7482;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_5 <= _GEN_4072;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_5 <= _GEN_7546;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_6 <= _GEN_4073;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_6 <= _GEN_7610;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_6_7 <= _GEN_4074;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_6_7 <= _GEN_7674;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_0 <= _GEN_4075;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_0 <= _GEN_7227;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_1 <= _GEN_4076;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_1 <= _GEN_7291;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_2 <= _GEN_4077;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_2 <= _GEN_7355;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_3 <= _GEN_4078;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_3 <= _GEN_7419;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_4 <= _GEN_4079;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_4 <= _GEN_7483;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_5 <= _GEN_4080;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_5 <= _GEN_7547;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_6 <= _GEN_4081;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_6 <= _GEN_7611;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_3_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_3_7_7 <= _GEN_4082;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_3_7_7 <= _GEN_7675;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_0 <= _GEN_4083;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_0 <= _GEN_7228;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_1 <= _GEN_4084;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_1 <= _GEN_7292;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_2 <= _GEN_4085;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_2 <= _GEN_7356;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_3 <= _GEN_4086;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_3 <= _GEN_7420;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_4 <= _GEN_4087;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_4 <= _GEN_7484;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_5 <= _GEN_4088;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_5 <= _GEN_7548;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_6 <= _GEN_4089;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_6 <= _GEN_7612;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_0_7 <= _GEN_4090;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_0_7 <= _GEN_7676;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_0 <= _GEN_4091;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_0 <= _GEN_7229;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_1 <= _GEN_4092;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_1 <= _GEN_7293;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_2 <= _GEN_4093;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_2 <= _GEN_7357;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_3 <= _GEN_4094;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_3 <= _GEN_7421;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_4 <= _GEN_4095;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_4 <= _GEN_7485;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_5 <= _GEN_4096;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_5 <= _GEN_7549;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_6 <= _GEN_4097;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_6 <= _GEN_7613;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_1_7 <= _GEN_4098;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_1_7 <= _GEN_7677;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_0 <= _GEN_4099;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_0 <= _GEN_7230;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_1 <= _GEN_4100;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_1 <= _GEN_7294;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_2 <= _GEN_4101;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_2 <= _GEN_7358;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_3 <= _GEN_4102;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_3 <= _GEN_7422;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_4 <= _GEN_4103;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_4 <= _GEN_7486;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_5 <= _GEN_4104;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_5 <= _GEN_7550;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_6 <= _GEN_4105;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_6 <= _GEN_7614;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_2_7 <= _GEN_4106;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_2_7 <= _GEN_7678;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_0 <= _GEN_4107;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_0 <= _GEN_7231;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_1 <= _GEN_4108;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_1 <= _GEN_7295;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_2 <= _GEN_4109;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_2 <= _GEN_7359;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_3 <= _GEN_4110;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_3 <= _GEN_7423;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_4 <= _GEN_4111;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_4 <= _GEN_7487;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_5 <= _GEN_4112;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_5 <= _GEN_7551;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_6 <= _GEN_4113;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_6 <= _GEN_7615;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_3_7 <= _GEN_4114;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_3_7 <= _GEN_7679;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_0 <= _GEN_4115;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_0 <= _GEN_7232;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_1 <= _GEN_4116;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_1 <= _GEN_7296;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_2 <= _GEN_4117;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_2 <= _GEN_7360;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_3 <= _GEN_4118;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_3 <= _GEN_7424;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_4 <= _GEN_4119;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_4 <= _GEN_7488;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_5 <= _GEN_4120;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_5 <= _GEN_7552;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_6 <= _GEN_4121;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_6 <= _GEN_7616;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_4_7 <= _GEN_4122;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_4_7 <= _GEN_7680;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_0 <= _GEN_4123;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_0 <= _GEN_7233;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_1 <= _GEN_4124;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_1 <= _GEN_7297;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_2 <= _GEN_4125;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_2 <= _GEN_7361;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_3 <= _GEN_4126;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_3 <= _GEN_7425;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_4 <= _GEN_4127;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_4 <= _GEN_7489;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_5 <= _GEN_4128;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_5 <= _GEN_7553;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_6 <= _GEN_4129;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_6 <= _GEN_7617;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_5_7 <= _GEN_4130;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_5_7 <= _GEN_7681;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_0 <= _GEN_4131;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_0 <= _GEN_7234;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_1 <= _GEN_4132;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_1 <= _GEN_7298;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_2 <= _GEN_4133;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_2 <= _GEN_7362;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_3 <= _GEN_4134;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_3 <= _GEN_7426;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_4 <= _GEN_4135;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_4 <= _GEN_7490;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_5 <= _GEN_4136;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_5 <= _GEN_7554;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_6 <= _GEN_4137;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_6 <= _GEN_7618;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_6_7 <= _GEN_4138;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_6_7 <= _GEN_7682;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_0 <= _GEN_4139;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_0 <= _GEN_7235;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_1 <= _GEN_4140;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_1 <= _GEN_7299;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_2 <= _GEN_4141;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_2 <= _GEN_7363;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_3 <= _GEN_4142;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_3 <= _GEN_7427;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_4 <= _GEN_4143;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_4 <= _GEN_7491;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_5 <= _GEN_4144;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_5 <= _GEN_7555;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_6 <= _GEN_4145;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_6 <= _GEN_7619;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_4_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_4_7_7 <= _GEN_4146;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_4_7_7 <= _GEN_7683;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_0 <= _GEN_4147;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_0 <= _GEN_7236;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_1 <= _GEN_4148;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_1 <= _GEN_7300;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_2 <= _GEN_4149;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_2 <= _GEN_7364;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_3 <= _GEN_4150;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_3 <= _GEN_7428;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_4 <= _GEN_4151;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_4 <= _GEN_7492;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_5 <= _GEN_4152;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_5 <= _GEN_7556;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_6 <= _GEN_4153;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_6 <= _GEN_7620;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_0_7 <= _GEN_4154;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_0_7 <= _GEN_7684;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_0 <= _GEN_4155;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_0 <= _GEN_7237;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_1 <= _GEN_4156;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_1 <= _GEN_7301;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_2 <= _GEN_4157;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_2 <= _GEN_7365;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_3 <= _GEN_4158;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_3 <= _GEN_7429;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_4 <= _GEN_4159;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_4 <= _GEN_7493;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_5 <= _GEN_4160;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_5 <= _GEN_7557;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_6 <= _GEN_4161;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_6 <= _GEN_7621;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_1_7 <= _GEN_4162;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_1_7 <= _GEN_7685;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_0 <= _GEN_4163;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_0 <= _GEN_7238;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_1 <= _GEN_4164;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_1 <= _GEN_7302;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_2 <= _GEN_4165;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_2 <= _GEN_7366;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_3 <= _GEN_4166;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_3 <= _GEN_7430;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_4 <= _GEN_4167;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_4 <= _GEN_7494;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_5 <= _GEN_4168;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_5 <= _GEN_7558;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_6 <= _GEN_4169;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_6 <= _GEN_7622;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_2_7 <= _GEN_4170;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_2_7 <= _GEN_7686;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_0 <= _GEN_4171;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_0 <= _GEN_7239;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_1 <= _GEN_4172;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_1 <= _GEN_7303;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_2 <= _GEN_4173;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_2 <= _GEN_7367;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_3 <= _GEN_4174;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_3 <= _GEN_7431;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_4 <= _GEN_4175;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_4 <= _GEN_7495;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_5 <= _GEN_4176;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_5 <= _GEN_7559;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_6 <= _GEN_4177;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_6 <= _GEN_7623;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_3_7 <= _GEN_4178;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_3_7 <= _GEN_7687;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_0 <= _GEN_4179;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_0 <= _GEN_7240;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_1 <= _GEN_4180;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_1 <= _GEN_7304;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_2 <= _GEN_4181;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_2 <= _GEN_7368;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_3 <= _GEN_4182;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_3 <= _GEN_7432;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_4 <= _GEN_4183;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_4 <= _GEN_7496;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_5 <= _GEN_4184;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_5 <= _GEN_7560;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_6 <= _GEN_4185;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_6 <= _GEN_7624;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_4_7 <= _GEN_4186;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_4_7 <= _GEN_7688;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_0 <= _GEN_4187;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_0 <= _GEN_7241;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_1 <= _GEN_4188;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_1 <= _GEN_7305;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_2 <= _GEN_4189;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_2 <= _GEN_7369;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_3 <= _GEN_4190;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_3 <= _GEN_7433;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_4 <= _GEN_4191;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_4 <= _GEN_7497;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_5 <= _GEN_4192;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_5 <= _GEN_7561;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_6 <= _GEN_4193;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_6 <= _GEN_7625;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_5_7 <= _GEN_4194;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_5_7 <= _GEN_7689;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_0 <= _GEN_4195;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_0 <= _GEN_7242;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_1 <= _GEN_4196;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_1 <= _GEN_7306;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_2 <= _GEN_4197;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_2 <= _GEN_7370;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_3 <= _GEN_4198;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_3 <= _GEN_7434;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_4 <= _GEN_4199;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_4 <= _GEN_7498;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_5 <= _GEN_4200;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_5 <= _GEN_7562;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_6 <= _GEN_4201;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_6 <= _GEN_7626;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_6_7 <= _GEN_4202;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_6_7 <= _GEN_7690;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_0 <= _GEN_4203;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_0 <= _GEN_7243;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_1 <= _GEN_4204;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_1 <= _GEN_7307;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_2 <= _GEN_4205;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_2 <= _GEN_7371;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_3 <= _GEN_4206;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_3 <= _GEN_7435;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_4 <= _GEN_4207;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_4 <= _GEN_7499;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_5 <= _GEN_4208;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_5 <= _GEN_7563;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_6 <= _GEN_4209;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_6 <= _GEN_7627;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_5_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_5_7_7 <= _GEN_4210;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_5_7_7 <= _GEN_7691;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_0 <= _GEN_4211;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_0 <= _GEN_7244;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_1 <= _GEN_4212;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_1 <= _GEN_7308;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_2 <= _GEN_4213;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_2 <= _GEN_7372;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_3 <= _GEN_4214;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_3 <= _GEN_7436;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_4 <= _GEN_4215;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_4 <= _GEN_7500;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_5 <= _GEN_4216;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_5 <= _GEN_7564;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_6 <= _GEN_4217;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_6 <= _GEN_7628;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_0_7 <= _GEN_4218;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_0_7 <= _GEN_7692;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_0 <= _GEN_4219;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_0 <= _GEN_7245;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_1 <= _GEN_4220;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_1 <= _GEN_7309;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_2 <= _GEN_4221;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_2 <= _GEN_7373;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_3 <= _GEN_4222;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_3 <= _GEN_7437;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_4 <= _GEN_4223;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_4 <= _GEN_7501;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_5 <= _GEN_4224;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_5 <= _GEN_7565;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_6 <= _GEN_4225;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_6 <= _GEN_7629;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_1_7 <= _GEN_4226;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_1_7 <= _GEN_7693;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_0 <= _GEN_4227;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_0 <= _GEN_7246;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_1 <= _GEN_4228;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_1 <= _GEN_7310;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_2 <= _GEN_4229;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_2 <= _GEN_7374;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_3 <= _GEN_4230;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_3 <= _GEN_7438;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_4 <= _GEN_4231;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_4 <= _GEN_7502;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_5 <= _GEN_4232;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_5 <= _GEN_7566;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_6 <= _GEN_4233;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_6 <= _GEN_7630;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_2_7 <= _GEN_4234;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_2_7 <= _GEN_7694;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_0 <= _GEN_4235;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_0 <= _GEN_7247;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_1 <= _GEN_4236;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_1 <= _GEN_7311;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_2 <= _GEN_4237;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_2 <= _GEN_7375;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_3 <= _GEN_4238;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_3 <= _GEN_7439;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_4 <= _GEN_4239;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_4 <= _GEN_7503;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_5 <= _GEN_4240;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_5 <= _GEN_7567;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_6 <= _GEN_4241;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_6 <= _GEN_7631;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_3_7 <= _GEN_4242;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_3_7 <= _GEN_7695;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_0 <= _GEN_4243;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_0 <= _GEN_7248;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_1 <= _GEN_4244;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_1 <= _GEN_7312;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_2 <= _GEN_4245;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_2 <= _GEN_7376;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_3 <= _GEN_4246;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_3 <= _GEN_7440;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_4 <= _GEN_4247;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_4 <= _GEN_7504;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_5 <= _GEN_4248;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_5 <= _GEN_7568;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_6 <= _GEN_4249;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_6 <= _GEN_7632;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_4_7 <= _GEN_4250;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_4_7 <= _GEN_7696;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_0 <= _GEN_4251;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_0 <= _GEN_7249;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_1 <= _GEN_4252;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_1 <= _GEN_7313;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_2 <= _GEN_4253;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_2 <= _GEN_7377;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_3 <= _GEN_4254;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_3 <= _GEN_7441;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_4 <= _GEN_4255;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_4 <= _GEN_7505;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_5 <= _GEN_4256;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_5 <= _GEN_7569;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_6 <= _GEN_4257;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_6 <= _GEN_7633;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_5_7 <= _GEN_4258;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_5_7 <= _GEN_7697;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_0 <= _GEN_4259;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_0 <= _GEN_7250;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_1 <= _GEN_4260;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_1 <= _GEN_7314;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_2 <= _GEN_4261;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_2 <= _GEN_7378;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_3 <= _GEN_4262;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_3 <= _GEN_7442;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_4 <= _GEN_4263;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_4 <= _GEN_7506;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_5 <= _GEN_4264;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_5 <= _GEN_7570;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_6 <= _GEN_4265;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_6 <= _GEN_7634;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_6_7 <= _GEN_4266;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_6_7 <= _GEN_7698;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_0 <= _GEN_4267;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_0 <= _GEN_7251;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_1 <= _GEN_4268;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_1 <= _GEN_7315;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_2 <= _GEN_4269;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_2 <= _GEN_7379;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_3 <= _GEN_4270;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_3 <= _GEN_7443;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_4 <= _GEN_4271;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_4 <= _GEN_7507;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_5 <= _GEN_4272;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_5 <= _GEN_7571;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_6 <= _GEN_4273;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_6 <= _GEN_7635;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_6_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_6_7_7 <= _GEN_4274;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_6_7_7 <= _GEN_7699;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_0 <= _GEN_4275;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_0 <= _GEN_7252;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_1 <= _GEN_4276;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_1 <= _GEN_7316;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_2 <= _GEN_4277;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_2 <= _GEN_7380;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_3 <= _GEN_4278;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_3 <= _GEN_7444;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_4 <= _GEN_4279;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_4 <= _GEN_7508;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_5 <= _GEN_4280;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_5 <= _GEN_7572;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_6 <= _GEN_4281;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_6 <= _GEN_7636;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_0_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_0_7 <= _GEN_4282;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_0_7 <= _GEN_7700;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_0 <= _GEN_4283;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_0 <= _GEN_7253;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_1 <= _GEN_4284;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_1 <= _GEN_7317;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_2 <= _GEN_4285;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_2 <= _GEN_7381;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_3 <= _GEN_4286;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_3 <= _GEN_7445;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_4 <= _GEN_4287;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_4 <= _GEN_7509;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_5 <= _GEN_4288;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_5 <= _GEN_7573;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_6 <= _GEN_4289;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_6 <= _GEN_7637;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_1_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_1_7 <= _GEN_4290;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_1_7 <= _GEN_7701;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_0 <= _GEN_4291;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_0 <= _GEN_7254;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_1 <= _GEN_4292;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_1 <= _GEN_7318;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_2 <= _GEN_4293;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_2 <= _GEN_7382;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_3 <= _GEN_4294;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_3 <= _GEN_7446;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_4 <= _GEN_4295;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_4 <= _GEN_7510;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_5 <= _GEN_4296;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_5 <= _GEN_7574;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_6 <= _GEN_4297;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_6 <= _GEN_7638;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_2_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_2_7 <= _GEN_4298;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_2_7 <= _GEN_7702;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_0 <= _GEN_4299;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_0 <= _GEN_7255;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_1 <= _GEN_4300;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_1 <= _GEN_7319;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_2 <= _GEN_4301;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_2 <= _GEN_7383;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_3 <= _GEN_4302;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_3 <= _GEN_7447;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_4 <= _GEN_4303;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_4 <= _GEN_7511;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_5 <= _GEN_4304;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_5 <= _GEN_7575;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_6 <= _GEN_4305;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_6 <= _GEN_7639;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_3_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_3_7 <= _GEN_4306;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_3_7 <= _GEN_7703;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_0 <= _GEN_4307;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_0 <= _GEN_7256;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_1 <= _GEN_4308;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_1 <= _GEN_7320;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_2 <= _GEN_4309;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_2 <= _GEN_7384;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_3 <= _GEN_4310;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_3 <= _GEN_7448;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_4 <= _GEN_4311;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_4 <= _GEN_7512;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_5 <= _GEN_4312;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_5 <= _GEN_7576;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_6 <= _GEN_4313;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_6 <= _GEN_7640;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_4_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_4_7 <= _GEN_4314;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_4_7 <= _GEN_7704;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_0 <= _GEN_4315;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_0 <= _GEN_7257;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_1 <= _GEN_4316;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_1 <= _GEN_7321;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_2 <= _GEN_4317;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_2 <= _GEN_7385;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_3 <= _GEN_4318;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_3 <= _GEN_7449;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_4 <= _GEN_4319;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_4 <= _GEN_7513;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_5 <= _GEN_4320;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_5 <= _GEN_7577;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_6 <= _GEN_4321;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_6 <= _GEN_7641;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_5_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_5_7 <= _GEN_4322;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_5_7 <= _GEN_7705;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_0 <= _GEN_4323;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_0 <= _GEN_7258;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_1 <= _GEN_4324;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_1 <= _GEN_7322;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_2 <= _GEN_4325;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_2 <= _GEN_7386;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_3 <= _GEN_4326;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_3 <= _GEN_7450;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_4 <= _GEN_4327;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_4 <= _GEN_7514;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_5 <= _GEN_4328;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_5 <= _GEN_7578;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_6 <= _GEN_4329;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_6 <= _GEN_7642;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_6_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_6_7 <= _GEN_4330;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_6_7 <= _GEN_7706;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_0 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_0 <= _GEN_4331;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_0 <= _GEN_7259;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_1 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_1 <= _GEN_4332;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_1 <= _GEN_7323;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_2 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_2 <= _GEN_4333;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_2 <= _GEN_7387;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_3 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_3 <= _GEN_4334;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_3 <= _GEN_7451;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_4 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_4 <= _GEN_4335;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_4 <= _GEN_7515;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_5 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_5 <= _GEN_4336;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_5 <= _GEN_7579;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_6 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_6 <= _GEN_4337;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_6 <= _GEN_7643;
      end
    end
    if (reset) begin // @[Cache.scala 53:25]
      CacheMem_7_7_7 <= 32'h0; // @[Cache.scala 53:25]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          CacheMem_7_7_7 <= _GEN_4338;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        CacheMem_7_7_7 <= _GEN_7707;
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_0 <= _GEN_7004;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_1 <= _GEN_7005;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_2 <= _GEN_7006;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_3 <= _GEN_7007;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_4 <= _GEN_7008;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_5 <= _GEN_7009;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_6 <= _GEN_7010;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_0_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_0_7 <= _GEN_7011;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_0 <= _GEN_7012;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_1 <= _GEN_7013;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_2 <= _GEN_7014;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_3 <= _GEN_7015;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_4 <= _GEN_7016;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_5 <= _GEN_7017;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_6 <= _GEN_7018;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_1_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_1_7 <= _GEN_7019;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_0 <= _GEN_7020;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_1 <= _GEN_7021;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_2 <= _GEN_7022;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_3 <= _GEN_7023;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_4 <= _GEN_7024;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_5 <= _GEN_7025;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_6 <= _GEN_7026;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_2_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_2_7 <= _GEN_7027;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_0 <= _GEN_7028;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_1 <= _GEN_7029;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_2 <= _GEN_7030;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_3 <= _GEN_7031;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_4 <= _GEN_7032;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_5 <= _GEN_7033;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_6 <= _GEN_7034;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_3_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_3_7 <= _GEN_7035;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_0 <= _GEN_7036;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_1 <= _GEN_7037;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_2 <= _GEN_7038;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_3 <= _GEN_7039;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_4 <= _GEN_7040;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_5 <= _GEN_7041;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_6 <= _GEN_7042;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_4_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_4_7 <= _GEN_7043;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_0 <= _GEN_7044;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_1 <= _GEN_7045;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_2 <= _GEN_7046;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_3 <= _GEN_7047;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_4 <= _GEN_7048;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_5 <= _GEN_7049;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_6 <= _GEN_7050;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_5_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_5_7 <= _GEN_7051;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_0 <= _GEN_7052;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_1 <= _GEN_7053;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_2 <= _GEN_7054;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_3 <= _GEN_7055;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_4 <= _GEN_7056;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_5 <= _GEN_7057;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_6 <= _GEN_7058;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_6_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_6_7 <= _GEN_7059;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_0 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_0 <= _GEN_7060;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_1 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_1 <= _GEN_7061;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_2 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_2 <= _GEN_7062;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_3 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_3 <= _GEN_7063;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_4 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_4 <= _GEN_7064;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_5 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_5 <= _GEN_7065;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_6 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_6 <= _GEN_7066;
        end
      end
    end
    if (reset) begin // @[Cache.scala 56:27]
      cache_tags_7_7 <= 6'h0; // @[Cache.scala 56:27]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          cache_tags_7_7 <= _GEN_7067;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_0 <= _GEN_7068;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_1 <= _GEN_7069;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_2 <= _GEN_7070;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_3 <= _GEN_7071;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_4 <= _GEN_7072;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_5 <= _GEN_7073;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_6 <= _GEN_7074;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_0_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_0_7 <= _GEN_7075;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_0 <= _GEN_7076;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_1 <= _GEN_7077;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_2 <= _GEN_7078;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_3 <= _GEN_7079;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_4 <= _GEN_7080;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_5 <= _GEN_7081;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_6 <= _GEN_7082;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_1_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_1_7 <= _GEN_7083;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_0 <= _GEN_7084;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_1 <= _GEN_7085;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_2 <= _GEN_7086;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_3 <= _GEN_7087;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_4 <= _GEN_7088;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_5 <= _GEN_7089;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_6 <= _GEN_7090;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_2_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_2_7 <= _GEN_7091;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_0 <= _GEN_7092;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_1 <= _GEN_7093;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_2 <= _GEN_7094;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_3 <= _GEN_7095;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_4 <= _GEN_7096;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_5 <= _GEN_7097;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_6 <= _GEN_7098;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_3_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_3_7 <= _GEN_7099;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_0 <= _GEN_7100;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_1 <= _GEN_7101;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_2 <= _GEN_7102;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_3 <= _GEN_7103;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_4 <= _GEN_7104;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_5 <= _GEN_7105;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_6 <= _GEN_7106;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_4_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_4_7 <= _GEN_7107;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_0 <= _GEN_7108;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_1 <= _GEN_7109;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_2 <= _GEN_7110;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_3 <= _GEN_7111;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_4 <= _GEN_7112;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_5 <= _GEN_7113;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_6 <= _GEN_7114;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_5_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_5_7 <= _GEN_7115;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_0 <= _GEN_7116;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_1 <= _GEN_7117;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_2 <= _GEN_7118;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_3 <= _GEN_7119;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_4 <= _GEN_7120;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_5 <= _GEN_7121;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_6 <= _GEN_7122;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_6_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_6_7 <= _GEN_7123;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_0 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_0 <= _GEN_7124;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_1 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_1 <= _GEN_7125;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_2 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_2 <= _GEN_7126;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_3 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_3 <= _GEN_7127;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_4 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_4 <= _GEN_7128;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_5 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_5 <= _GEN_7129;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_6 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_6 <= _GEN_7130;
        end
      end
    end
    if (reset) begin // @[Cache.scala 57:22]
      valid_7_7 <= 1'h0; // @[Cache.scala 57:22]
    end else if (!(_T_27)) begin // @[Cache.scala 126:21]
      if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
        if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
          valid_7_7 <= _GEN_7131;
        end
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_0 <= _GEN_4339;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_0 <= _GEN_7132;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_1 <= _GEN_4340;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_1 <= _GEN_7133;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_2 <= _GEN_4341;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_2 <= _GEN_7134;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_3 <= _GEN_4342;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_3 <= _GEN_7135;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_4 <= _GEN_4343;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_4 <= _GEN_7136;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_5 <= _GEN_4344;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_5 <= _GEN_7137;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_6 <= _GEN_4345;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_6 <= _GEN_7138;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_0_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_0_7 <= _GEN_4346;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_0_7 <= _GEN_7139;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_0 <= _GEN_4347;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_0 <= _GEN_7140;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_1 <= _GEN_4348;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_1 <= _GEN_7141;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_2 <= _GEN_4349;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_2 <= _GEN_7142;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_3 <= _GEN_4350;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_3 <= _GEN_7143;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_4 <= _GEN_4351;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_4 <= _GEN_7144;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_5 <= _GEN_4352;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_5 <= _GEN_7145;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_6 <= _GEN_4353;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_6 <= _GEN_7146;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_1_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_1_7 <= _GEN_4354;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_1_7 <= _GEN_7147;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_0 <= _GEN_4355;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_0 <= _GEN_7148;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_1 <= _GEN_4356;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_1 <= _GEN_7149;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_2 <= _GEN_4357;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_2 <= _GEN_7150;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_3 <= _GEN_4358;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_3 <= _GEN_7151;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_4 <= _GEN_4359;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_4 <= _GEN_7152;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_5 <= _GEN_4360;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_5 <= _GEN_7153;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_6 <= _GEN_4361;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_6 <= _GEN_7154;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_2_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_2_7 <= _GEN_4362;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_2_7 <= _GEN_7155;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_0 <= _GEN_4363;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_0 <= _GEN_7156;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_1 <= _GEN_4364;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_1 <= _GEN_7157;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_2 <= _GEN_4365;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_2 <= _GEN_7158;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_3 <= _GEN_4366;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_3 <= _GEN_7159;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_4 <= _GEN_4367;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_4 <= _GEN_7160;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_5 <= _GEN_4368;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_5 <= _GEN_7161;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_6 <= _GEN_4369;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_6 <= _GEN_7162;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_3_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_3_7 <= _GEN_4370;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_3_7 <= _GEN_7163;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_0 <= _GEN_4371;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_0 <= _GEN_7164;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_1 <= _GEN_4372;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_1 <= _GEN_7165;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_2 <= _GEN_4373;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_2 <= _GEN_7166;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_3 <= _GEN_4374;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_3 <= _GEN_7167;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_4 <= _GEN_4375;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_4 <= _GEN_7168;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_5 <= _GEN_4376;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_5 <= _GEN_7169;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_6 <= _GEN_4377;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_6 <= _GEN_7170;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_4_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_4_7 <= _GEN_4378;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_4_7 <= _GEN_7171;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_0 <= _GEN_4379;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_0 <= _GEN_7172;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_1 <= _GEN_4380;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_1 <= _GEN_7173;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_2 <= _GEN_4381;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_2 <= _GEN_7174;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_3 <= _GEN_4382;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_3 <= _GEN_7175;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_4 <= _GEN_4383;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_4 <= _GEN_7176;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_5 <= _GEN_4384;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_5 <= _GEN_7177;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_6 <= _GEN_4385;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_6 <= _GEN_7178;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_5_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_5_7 <= _GEN_4386;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_5_7 <= _GEN_7179;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_0 <= _GEN_4387;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_0 <= _GEN_7180;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_1 <= _GEN_4388;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_1 <= _GEN_7181;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_2 <= _GEN_4389;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_2 <= _GEN_7182;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_3 <= _GEN_4390;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_3 <= _GEN_7183;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_4 <= _GEN_4391;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_4 <= _GEN_7184;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_5 <= _GEN_4392;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_5 <= _GEN_7185;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_6 <= _GEN_4393;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_6 <= _GEN_7186;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_6_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_6_7 <= _GEN_4394;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_6_7 <= _GEN_7187;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_0 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_0 <= _GEN_4395;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_0 <= _GEN_7188;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_1 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_1 <= _GEN_4396;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_1 <= _GEN_7189;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_2 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_2 <= _GEN_4397;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_2 <= _GEN_7190;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_3 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_3 <= _GEN_4398;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_3 <= _GEN_7191;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_4 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_4 <= _GEN_4399;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_4 <= _GEN_7192;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_5 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_5 <= _GEN_4400;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_5 <= _GEN_7193;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_6 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_6 <= _GEN_4401;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_6 <= _GEN_7194;
      end
    end
    if (reset) begin // @[Cache.scala 58:22]
      dirty_7_7 <= 1'h0; // @[Cache.scala 58:22]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          dirty_7_7 <= _GEN_4402;
        end
      end
    end else if (!(2'h1 == cacheState)) begin // @[Cache.scala 126:21]
      if (!(2'h2 == cacheState)) begin // @[Cache.scala 126:21]
        dirty_7_7 <= _GEN_7195;
      end
    end
    if (reset) begin // @[Cache.scala 70:32]
      mem_rd_set_addr <= 3'h0; // @[Cache.scala 70:32]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_rd_set_addr <= set_addr; // @[Cache.scala 158:27]
        end
      end
    end
    if (reset) begin // @[Cache.scala 71:32]
      mem_rd_tag_addr <= 6'h0; // @[Cache.scala 71:32]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_rd_tag_addr <= tag_addr; // @[Cache.scala 157:27]
        end
      end
    end
    if (reset) begin // @[Cache.scala 73:28]
      mem_wr_addr <= 9'h0; // @[Cache.scala 73:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_addr <= _GEN_5687;
        end
      end
    end
    if (reset) begin // @[Cache.scala 96:27]
      cacheState <= 2'h0; // @[Cache.scala 96:27]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (cache_Hit) begin // @[Cache.scala 128:22]
        if (!(io_r_req)) begin // @[Cache.scala 129:34]
          cacheState <= _GEN_4403;
        end
      end else if (_T) begin // @[Cache.scala 149:34]
        cacheState <= _GEN_5686;
      end
    end else if (2'h1 == cacheState) begin // @[Cache.scala 126:21]
      if (io_cacheAXI_gnt) begin // @[Cache.scala 163:39]
        cacheState <= 2'h2; // @[Cache.scala 164:20]
      end
    end else if (2'h2 == cacheState) begin // @[Cache.scala 126:21]
      cacheState <= _GEN_6298;
    end else begin
      cacheState <= _GEN_7003;
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_0 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h0 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_0 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_1 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h1 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_1 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_2 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h2 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_2 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_3 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h3 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_3 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_4 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h4 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_4 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_5 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h5 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_5 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_6 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h6 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_6 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 103:30]
      FIFO_Choice_7 <= 32'h0; // @[Cache.scala 103:30]
    end else if (!(2'h0 == cacheState)) begin // @[Cache.scala 104:23]
      if (2'h3 == cacheState) begin // @[Cache.scala 104:23]
        if (3'h7 == set_addr) begin // @[Cache.scala 109:31]
          FIFO_Choice_7 <= _FIFO_Choice_set_addr_1; // @[Cache.scala 109:31]
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_0 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_0 <= _GEN_5688;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_1 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_1 <= _GEN_5689;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_2 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_2 <= _GEN_5690;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_3 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_3 <= _GEN_5691;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_4 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_4 <= _GEN_5692;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_5 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_5 <= _GEN_5693;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_6 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_6 <= _GEN_5694;
        end
      end
    end
    if (reset) begin // @[Cache.scala 124:28]
      mem_wr_line_7 <= 32'h0; // @[Cache.scala 124:28]
    end else if (_T_27) begin // @[Cache.scala 126:21]
      if (!(cache_Hit)) begin // @[Cache.scala 128:22]
        if (_T) begin // @[Cache.scala 149:34]
          mem_wr_line_7 <= _GEN_5695;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  CacheMem_0_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  CacheMem_0_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  CacheMem_0_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  CacheMem_0_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  CacheMem_0_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  CacheMem_0_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  CacheMem_0_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  CacheMem_0_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  CacheMem_0_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  CacheMem_0_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  CacheMem_0_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  CacheMem_0_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  CacheMem_0_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  CacheMem_0_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  CacheMem_0_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  CacheMem_0_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  CacheMem_0_2_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  CacheMem_0_2_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  CacheMem_0_2_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  CacheMem_0_2_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  CacheMem_0_2_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  CacheMem_0_2_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  CacheMem_0_2_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  CacheMem_0_2_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  CacheMem_0_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  CacheMem_0_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  CacheMem_0_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  CacheMem_0_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  CacheMem_0_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  CacheMem_0_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  CacheMem_0_3_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  CacheMem_0_3_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  CacheMem_0_4_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  CacheMem_0_4_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  CacheMem_0_4_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  CacheMem_0_4_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  CacheMem_0_4_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  CacheMem_0_4_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  CacheMem_0_4_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  CacheMem_0_4_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  CacheMem_0_5_0 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  CacheMem_0_5_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  CacheMem_0_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  CacheMem_0_5_3 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  CacheMem_0_5_4 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  CacheMem_0_5_5 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  CacheMem_0_5_6 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  CacheMem_0_5_7 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  CacheMem_0_6_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  CacheMem_0_6_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  CacheMem_0_6_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  CacheMem_0_6_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  CacheMem_0_6_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  CacheMem_0_6_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  CacheMem_0_6_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  CacheMem_0_6_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  CacheMem_0_7_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  CacheMem_0_7_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  CacheMem_0_7_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  CacheMem_0_7_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  CacheMem_0_7_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  CacheMem_0_7_5 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  CacheMem_0_7_6 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  CacheMem_0_7_7 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  CacheMem_1_0_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  CacheMem_1_0_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  CacheMem_1_0_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  CacheMem_1_0_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  CacheMem_1_0_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  CacheMem_1_0_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  CacheMem_1_0_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  CacheMem_1_0_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  CacheMem_1_1_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  CacheMem_1_1_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  CacheMem_1_1_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  CacheMem_1_1_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  CacheMem_1_1_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  CacheMem_1_1_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  CacheMem_1_1_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  CacheMem_1_1_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  CacheMem_1_2_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  CacheMem_1_2_1 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  CacheMem_1_2_2 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  CacheMem_1_2_3 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  CacheMem_1_2_4 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  CacheMem_1_2_5 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  CacheMem_1_2_6 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  CacheMem_1_2_7 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  CacheMem_1_3_0 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  CacheMem_1_3_1 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  CacheMem_1_3_2 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  CacheMem_1_3_3 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  CacheMem_1_3_4 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  CacheMem_1_3_5 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  CacheMem_1_3_6 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  CacheMem_1_3_7 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  CacheMem_1_4_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  CacheMem_1_4_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  CacheMem_1_4_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  CacheMem_1_4_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  CacheMem_1_4_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  CacheMem_1_4_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  CacheMem_1_4_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  CacheMem_1_4_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  CacheMem_1_5_0 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  CacheMem_1_5_1 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  CacheMem_1_5_2 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  CacheMem_1_5_3 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  CacheMem_1_5_4 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  CacheMem_1_5_5 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  CacheMem_1_5_6 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  CacheMem_1_5_7 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  CacheMem_1_6_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  CacheMem_1_6_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  CacheMem_1_6_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  CacheMem_1_6_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  CacheMem_1_6_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  CacheMem_1_6_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  CacheMem_1_6_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  CacheMem_1_6_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  CacheMem_1_7_0 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  CacheMem_1_7_1 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  CacheMem_1_7_2 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  CacheMem_1_7_3 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  CacheMem_1_7_4 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  CacheMem_1_7_5 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  CacheMem_1_7_6 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  CacheMem_1_7_7 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  CacheMem_2_0_0 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  CacheMem_2_0_1 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  CacheMem_2_0_2 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  CacheMem_2_0_3 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  CacheMem_2_0_4 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  CacheMem_2_0_5 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  CacheMem_2_0_6 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  CacheMem_2_0_7 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  CacheMem_2_1_0 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  CacheMem_2_1_1 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  CacheMem_2_1_2 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  CacheMem_2_1_3 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  CacheMem_2_1_4 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  CacheMem_2_1_5 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  CacheMem_2_1_6 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  CacheMem_2_1_7 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  CacheMem_2_2_0 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  CacheMem_2_2_1 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  CacheMem_2_2_2 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  CacheMem_2_2_3 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  CacheMem_2_2_4 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  CacheMem_2_2_5 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  CacheMem_2_2_6 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  CacheMem_2_2_7 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  CacheMem_2_3_0 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  CacheMem_2_3_1 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  CacheMem_2_3_2 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  CacheMem_2_3_3 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  CacheMem_2_3_4 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  CacheMem_2_3_5 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  CacheMem_2_3_6 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  CacheMem_2_3_7 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  CacheMem_2_4_0 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  CacheMem_2_4_1 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  CacheMem_2_4_2 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  CacheMem_2_4_3 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  CacheMem_2_4_4 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  CacheMem_2_4_5 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  CacheMem_2_4_6 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  CacheMem_2_4_7 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  CacheMem_2_5_0 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  CacheMem_2_5_1 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  CacheMem_2_5_2 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  CacheMem_2_5_3 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  CacheMem_2_5_4 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  CacheMem_2_5_5 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  CacheMem_2_5_6 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  CacheMem_2_5_7 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  CacheMem_2_6_0 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  CacheMem_2_6_1 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  CacheMem_2_6_2 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  CacheMem_2_6_3 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  CacheMem_2_6_4 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  CacheMem_2_6_5 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  CacheMem_2_6_6 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  CacheMem_2_6_7 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  CacheMem_2_7_0 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  CacheMem_2_7_1 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  CacheMem_2_7_2 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  CacheMem_2_7_3 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  CacheMem_2_7_4 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  CacheMem_2_7_5 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  CacheMem_2_7_6 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  CacheMem_2_7_7 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  CacheMem_3_0_0 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  CacheMem_3_0_1 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  CacheMem_3_0_2 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  CacheMem_3_0_3 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  CacheMem_3_0_4 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  CacheMem_3_0_5 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  CacheMem_3_0_6 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  CacheMem_3_0_7 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  CacheMem_3_1_0 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  CacheMem_3_1_1 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  CacheMem_3_1_2 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  CacheMem_3_1_3 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  CacheMem_3_1_4 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  CacheMem_3_1_5 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  CacheMem_3_1_6 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  CacheMem_3_1_7 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  CacheMem_3_2_0 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  CacheMem_3_2_1 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  CacheMem_3_2_2 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  CacheMem_3_2_3 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  CacheMem_3_2_4 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  CacheMem_3_2_5 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  CacheMem_3_2_6 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  CacheMem_3_2_7 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  CacheMem_3_3_0 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  CacheMem_3_3_1 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  CacheMem_3_3_2 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  CacheMem_3_3_3 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  CacheMem_3_3_4 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  CacheMem_3_3_5 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  CacheMem_3_3_6 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  CacheMem_3_3_7 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  CacheMem_3_4_0 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  CacheMem_3_4_1 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  CacheMem_3_4_2 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  CacheMem_3_4_3 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  CacheMem_3_4_4 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  CacheMem_3_4_5 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  CacheMem_3_4_6 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  CacheMem_3_4_7 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  CacheMem_3_5_0 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  CacheMem_3_5_1 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  CacheMem_3_5_2 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  CacheMem_3_5_3 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  CacheMem_3_5_4 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  CacheMem_3_5_5 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  CacheMem_3_5_6 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  CacheMem_3_5_7 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  CacheMem_3_6_0 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  CacheMem_3_6_1 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  CacheMem_3_6_2 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  CacheMem_3_6_3 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  CacheMem_3_6_4 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  CacheMem_3_6_5 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  CacheMem_3_6_6 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  CacheMem_3_6_7 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  CacheMem_3_7_0 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  CacheMem_3_7_1 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  CacheMem_3_7_2 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  CacheMem_3_7_3 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  CacheMem_3_7_4 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  CacheMem_3_7_5 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  CacheMem_3_7_6 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  CacheMem_3_7_7 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  CacheMem_4_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  CacheMem_4_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  CacheMem_4_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  CacheMem_4_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  CacheMem_4_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  CacheMem_4_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  CacheMem_4_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  CacheMem_4_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  CacheMem_4_1_0 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  CacheMem_4_1_1 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  CacheMem_4_1_2 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  CacheMem_4_1_3 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  CacheMem_4_1_4 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  CacheMem_4_1_5 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  CacheMem_4_1_6 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  CacheMem_4_1_7 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  CacheMem_4_2_0 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  CacheMem_4_2_1 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  CacheMem_4_2_2 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  CacheMem_4_2_3 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  CacheMem_4_2_4 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  CacheMem_4_2_5 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  CacheMem_4_2_6 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  CacheMem_4_2_7 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  CacheMem_4_3_0 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  CacheMem_4_3_1 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  CacheMem_4_3_2 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  CacheMem_4_3_3 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  CacheMem_4_3_4 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  CacheMem_4_3_5 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  CacheMem_4_3_6 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  CacheMem_4_3_7 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  CacheMem_4_4_0 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  CacheMem_4_4_1 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  CacheMem_4_4_2 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  CacheMem_4_4_3 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  CacheMem_4_4_4 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  CacheMem_4_4_5 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  CacheMem_4_4_6 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  CacheMem_4_4_7 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  CacheMem_4_5_0 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  CacheMem_4_5_1 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  CacheMem_4_5_2 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  CacheMem_4_5_3 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  CacheMem_4_5_4 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  CacheMem_4_5_5 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  CacheMem_4_5_6 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  CacheMem_4_5_7 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  CacheMem_4_6_0 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  CacheMem_4_6_1 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  CacheMem_4_6_2 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  CacheMem_4_6_3 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  CacheMem_4_6_4 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  CacheMem_4_6_5 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  CacheMem_4_6_6 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  CacheMem_4_6_7 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  CacheMem_4_7_0 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  CacheMem_4_7_1 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  CacheMem_4_7_2 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  CacheMem_4_7_3 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  CacheMem_4_7_4 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  CacheMem_4_7_5 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  CacheMem_4_7_6 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  CacheMem_4_7_7 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  CacheMem_5_0_0 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  CacheMem_5_0_1 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  CacheMem_5_0_2 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  CacheMem_5_0_3 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  CacheMem_5_0_4 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  CacheMem_5_0_5 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  CacheMem_5_0_6 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  CacheMem_5_0_7 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  CacheMem_5_1_0 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  CacheMem_5_1_1 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  CacheMem_5_1_2 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  CacheMem_5_1_3 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  CacheMem_5_1_4 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  CacheMem_5_1_5 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  CacheMem_5_1_6 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  CacheMem_5_1_7 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  CacheMem_5_2_0 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  CacheMem_5_2_1 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  CacheMem_5_2_2 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  CacheMem_5_2_3 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  CacheMem_5_2_4 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  CacheMem_5_2_5 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  CacheMem_5_2_6 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  CacheMem_5_2_7 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  CacheMem_5_3_0 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  CacheMem_5_3_1 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  CacheMem_5_3_2 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  CacheMem_5_3_3 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  CacheMem_5_3_4 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  CacheMem_5_3_5 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  CacheMem_5_3_6 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  CacheMem_5_3_7 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  CacheMem_5_4_0 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  CacheMem_5_4_1 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  CacheMem_5_4_2 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  CacheMem_5_4_3 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  CacheMem_5_4_4 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  CacheMem_5_4_5 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  CacheMem_5_4_6 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  CacheMem_5_4_7 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  CacheMem_5_5_0 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  CacheMem_5_5_1 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  CacheMem_5_5_2 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  CacheMem_5_5_3 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  CacheMem_5_5_4 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  CacheMem_5_5_5 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  CacheMem_5_5_6 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  CacheMem_5_5_7 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  CacheMem_5_6_0 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  CacheMem_5_6_1 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  CacheMem_5_6_2 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  CacheMem_5_6_3 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  CacheMem_5_6_4 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  CacheMem_5_6_5 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  CacheMem_5_6_6 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  CacheMem_5_6_7 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  CacheMem_5_7_0 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  CacheMem_5_7_1 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  CacheMem_5_7_2 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  CacheMem_5_7_3 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  CacheMem_5_7_4 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  CacheMem_5_7_5 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  CacheMem_5_7_6 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  CacheMem_5_7_7 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  CacheMem_6_0_0 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  CacheMem_6_0_1 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  CacheMem_6_0_2 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  CacheMem_6_0_3 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  CacheMem_6_0_4 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  CacheMem_6_0_5 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  CacheMem_6_0_6 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  CacheMem_6_0_7 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  CacheMem_6_1_0 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  CacheMem_6_1_1 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  CacheMem_6_1_2 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  CacheMem_6_1_3 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  CacheMem_6_1_4 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  CacheMem_6_1_5 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  CacheMem_6_1_6 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  CacheMem_6_1_7 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  CacheMem_6_2_0 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  CacheMem_6_2_1 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  CacheMem_6_2_2 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  CacheMem_6_2_3 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  CacheMem_6_2_4 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  CacheMem_6_2_5 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  CacheMem_6_2_6 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  CacheMem_6_2_7 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  CacheMem_6_3_0 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  CacheMem_6_3_1 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  CacheMem_6_3_2 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  CacheMem_6_3_3 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  CacheMem_6_3_4 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  CacheMem_6_3_5 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  CacheMem_6_3_6 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  CacheMem_6_3_7 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  CacheMem_6_4_0 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  CacheMem_6_4_1 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  CacheMem_6_4_2 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  CacheMem_6_4_3 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  CacheMem_6_4_4 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  CacheMem_6_4_5 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  CacheMem_6_4_6 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  CacheMem_6_4_7 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  CacheMem_6_5_0 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  CacheMem_6_5_1 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  CacheMem_6_5_2 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  CacheMem_6_5_3 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  CacheMem_6_5_4 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  CacheMem_6_5_5 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  CacheMem_6_5_6 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  CacheMem_6_5_7 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  CacheMem_6_6_0 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  CacheMem_6_6_1 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  CacheMem_6_6_2 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  CacheMem_6_6_3 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  CacheMem_6_6_4 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  CacheMem_6_6_5 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  CacheMem_6_6_6 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  CacheMem_6_6_7 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  CacheMem_6_7_0 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  CacheMem_6_7_1 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  CacheMem_6_7_2 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  CacheMem_6_7_3 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  CacheMem_6_7_4 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  CacheMem_6_7_5 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  CacheMem_6_7_6 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  CacheMem_6_7_7 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  CacheMem_7_0_0 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  CacheMem_7_0_1 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  CacheMem_7_0_2 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  CacheMem_7_0_3 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  CacheMem_7_0_4 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  CacheMem_7_0_5 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  CacheMem_7_0_6 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  CacheMem_7_0_7 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  CacheMem_7_1_0 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  CacheMem_7_1_1 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  CacheMem_7_1_2 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  CacheMem_7_1_3 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  CacheMem_7_1_4 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  CacheMem_7_1_5 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  CacheMem_7_1_6 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  CacheMem_7_1_7 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  CacheMem_7_2_0 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  CacheMem_7_2_1 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  CacheMem_7_2_2 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  CacheMem_7_2_3 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  CacheMem_7_2_4 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  CacheMem_7_2_5 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  CacheMem_7_2_6 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  CacheMem_7_2_7 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  CacheMem_7_3_0 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  CacheMem_7_3_1 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  CacheMem_7_3_2 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  CacheMem_7_3_3 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  CacheMem_7_3_4 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  CacheMem_7_3_5 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  CacheMem_7_3_6 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  CacheMem_7_3_7 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  CacheMem_7_4_0 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  CacheMem_7_4_1 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  CacheMem_7_4_2 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  CacheMem_7_4_3 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  CacheMem_7_4_4 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  CacheMem_7_4_5 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  CacheMem_7_4_6 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  CacheMem_7_4_7 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  CacheMem_7_5_0 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  CacheMem_7_5_1 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  CacheMem_7_5_2 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  CacheMem_7_5_3 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  CacheMem_7_5_4 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  CacheMem_7_5_5 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  CacheMem_7_5_6 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  CacheMem_7_5_7 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  CacheMem_7_6_0 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  CacheMem_7_6_1 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  CacheMem_7_6_2 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  CacheMem_7_6_3 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  CacheMem_7_6_4 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  CacheMem_7_6_5 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  CacheMem_7_6_6 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  CacheMem_7_6_7 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  CacheMem_7_7_0 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  CacheMem_7_7_1 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  CacheMem_7_7_2 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  CacheMem_7_7_3 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  CacheMem_7_7_4 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  CacheMem_7_7_5 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  CacheMem_7_7_6 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  CacheMem_7_7_7 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  cache_tags_0_0 = _RAND_512[5:0];
  _RAND_513 = {1{`RANDOM}};
  cache_tags_0_1 = _RAND_513[5:0];
  _RAND_514 = {1{`RANDOM}};
  cache_tags_0_2 = _RAND_514[5:0];
  _RAND_515 = {1{`RANDOM}};
  cache_tags_0_3 = _RAND_515[5:0];
  _RAND_516 = {1{`RANDOM}};
  cache_tags_0_4 = _RAND_516[5:0];
  _RAND_517 = {1{`RANDOM}};
  cache_tags_0_5 = _RAND_517[5:0];
  _RAND_518 = {1{`RANDOM}};
  cache_tags_0_6 = _RAND_518[5:0];
  _RAND_519 = {1{`RANDOM}};
  cache_tags_0_7 = _RAND_519[5:0];
  _RAND_520 = {1{`RANDOM}};
  cache_tags_1_0 = _RAND_520[5:0];
  _RAND_521 = {1{`RANDOM}};
  cache_tags_1_1 = _RAND_521[5:0];
  _RAND_522 = {1{`RANDOM}};
  cache_tags_1_2 = _RAND_522[5:0];
  _RAND_523 = {1{`RANDOM}};
  cache_tags_1_3 = _RAND_523[5:0];
  _RAND_524 = {1{`RANDOM}};
  cache_tags_1_4 = _RAND_524[5:0];
  _RAND_525 = {1{`RANDOM}};
  cache_tags_1_5 = _RAND_525[5:0];
  _RAND_526 = {1{`RANDOM}};
  cache_tags_1_6 = _RAND_526[5:0];
  _RAND_527 = {1{`RANDOM}};
  cache_tags_1_7 = _RAND_527[5:0];
  _RAND_528 = {1{`RANDOM}};
  cache_tags_2_0 = _RAND_528[5:0];
  _RAND_529 = {1{`RANDOM}};
  cache_tags_2_1 = _RAND_529[5:0];
  _RAND_530 = {1{`RANDOM}};
  cache_tags_2_2 = _RAND_530[5:0];
  _RAND_531 = {1{`RANDOM}};
  cache_tags_2_3 = _RAND_531[5:0];
  _RAND_532 = {1{`RANDOM}};
  cache_tags_2_4 = _RAND_532[5:0];
  _RAND_533 = {1{`RANDOM}};
  cache_tags_2_5 = _RAND_533[5:0];
  _RAND_534 = {1{`RANDOM}};
  cache_tags_2_6 = _RAND_534[5:0];
  _RAND_535 = {1{`RANDOM}};
  cache_tags_2_7 = _RAND_535[5:0];
  _RAND_536 = {1{`RANDOM}};
  cache_tags_3_0 = _RAND_536[5:0];
  _RAND_537 = {1{`RANDOM}};
  cache_tags_3_1 = _RAND_537[5:0];
  _RAND_538 = {1{`RANDOM}};
  cache_tags_3_2 = _RAND_538[5:0];
  _RAND_539 = {1{`RANDOM}};
  cache_tags_3_3 = _RAND_539[5:0];
  _RAND_540 = {1{`RANDOM}};
  cache_tags_3_4 = _RAND_540[5:0];
  _RAND_541 = {1{`RANDOM}};
  cache_tags_3_5 = _RAND_541[5:0];
  _RAND_542 = {1{`RANDOM}};
  cache_tags_3_6 = _RAND_542[5:0];
  _RAND_543 = {1{`RANDOM}};
  cache_tags_3_7 = _RAND_543[5:0];
  _RAND_544 = {1{`RANDOM}};
  cache_tags_4_0 = _RAND_544[5:0];
  _RAND_545 = {1{`RANDOM}};
  cache_tags_4_1 = _RAND_545[5:0];
  _RAND_546 = {1{`RANDOM}};
  cache_tags_4_2 = _RAND_546[5:0];
  _RAND_547 = {1{`RANDOM}};
  cache_tags_4_3 = _RAND_547[5:0];
  _RAND_548 = {1{`RANDOM}};
  cache_tags_4_4 = _RAND_548[5:0];
  _RAND_549 = {1{`RANDOM}};
  cache_tags_4_5 = _RAND_549[5:0];
  _RAND_550 = {1{`RANDOM}};
  cache_tags_4_6 = _RAND_550[5:0];
  _RAND_551 = {1{`RANDOM}};
  cache_tags_4_7 = _RAND_551[5:0];
  _RAND_552 = {1{`RANDOM}};
  cache_tags_5_0 = _RAND_552[5:0];
  _RAND_553 = {1{`RANDOM}};
  cache_tags_5_1 = _RAND_553[5:0];
  _RAND_554 = {1{`RANDOM}};
  cache_tags_5_2 = _RAND_554[5:0];
  _RAND_555 = {1{`RANDOM}};
  cache_tags_5_3 = _RAND_555[5:0];
  _RAND_556 = {1{`RANDOM}};
  cache_tags_5_4 = _RAND_556[5:0];
  _RAND_557 = {1{`RANDOM}};
  cache_tags_5_5 = _RAND_557[5:0];
  _RAND_558 = {1{`RANDOM}};
  cache_tags_5_6 = _RAND_558[5:0];
  _RAND_559 = {1{`RANDOM}};
  cache_tags_5_7 = _RAND_559[5:0];
  _RAND_560 = {1{`RANDOM}};
  cache_tags_6_0 = _RAND_560[5:0];
  _RAND_561 = {1{`RANDOM}};
  cache_tags_6_1 = _RAND_561[5:0];
  _RAND_562 = {1{`RANDOM}};
  cache_tags_6_2 = _RAND_562[5:0];
  _RAND_563 = {1{`RANDOM}};
  cache_tags_6_3 = _RAND_563[5:0];
  _RAND_564 = {1{`RANDOM}};
  cache_tags_6_4 = _RAND_564[5:0];
  _RAND_565 = {1{`RANDOM}};
  cache_tags_6_5 = _RAND_565[5:0];
  _RAND_566 = {1{`RANDOM}};
  cache_tags_6_6 = _RAND_566[5:0];
  _RAND_567 = {1{`RANDOM}};
  cache_tags_6_7 = _RAND_567[5:0];
  _RAND_568 = {1{`RANDOM}};
  cache_tags_7_0 = _RAND_568[5:0];
  _RAND_569 = {1{`RANDOM}};
  cache_tags_7_1 = _RAND_569[5:0];
  _RAND_570 = {1{`RANDOM}};
  cache_tags_7_2 = _RAND_570[5:0];
  _RAND_571 = {1{`RANDOM}};
  cache_tags_7_3 = _RAND_571[5:0];
  _RAND_572 = {1{`RANDOM}};
  cache_tags_7_4 = _RAND_572[5:0];
  _RAND_573 = {1{`RANDOM}};
  cache_tags_7_5 = _RAND_573[5:0];
  _RAND_574 = {1{`RANDOM}};
  cache_tags_7_6 = _RAND_574[5:0];
  _RAND_575 = {1{`RANDOM}};
  cache_tags_7_7 = _RAND_575[5:0];
  _RAND_576 = {1{`RANDOM}};
  valid_0_0 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_0_1 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_0_2 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_0_3 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_0_4 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_0_5 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_0_6 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_0_7 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_1_0 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_1_1 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_1_2 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_1_3 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_1_4 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_1_5 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_1_6 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_1_7 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_2_0 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_2_1 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_2_2 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_2_3 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_2_4 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_2_5 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_2_6 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_2_7 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_3_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_3_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_3_2 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_3_3 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_3_4 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_3_5 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_3_6 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_3_7 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_4_0 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_4_1 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_4_2 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_4_3 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_4_4 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_4_5 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_4_6 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_4_7 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_5_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_5_1 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_5_2 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_5_3 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_5_4 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_5_5 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_5_6 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_5_7 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_6_0 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_6_1 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_6_2 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_6_3 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_6_4 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_6_5 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_6_6 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_6_7 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_7_0 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_7_1 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_7_2 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_7_3 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_7_4 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_7_5 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_7_6 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_7_7 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  dirty_0_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  dirty_0_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  dirty_0_2 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  dirty_0_3 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  dirty_0_4 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  dirty_0_5 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  dirty_0_6 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  dirty_0_7 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  dirty_1_0 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  dirty_1_1 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  dirty_1_2 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  dirty_1_3 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  dirty_1_4 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  dirty_1_5 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  dirty_1_6 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  dirty_1_7 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  dirty_2_0 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  dirty_2_1 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  dirty_2_2 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  dirty_2_3 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  dirty_2_4 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  dirty_2_5 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  dirty_2_6 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  dirty_2_7 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  dirty_3_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  dirty_3_1 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  dirty_3_2 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  dirty_3_3 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  dirty_3_4 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  dirty_3_5 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  dirty_3_6 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  dirty_3_7 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  dirty_4_0 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  dirty_4_1 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  dirty_4_2 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  dirty_4_3 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  dirty_4_4 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  dirty_4_5 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  dirty_4_6 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  dirty_4_7 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  dirty_5_0 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  dirty_5_1 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  dirty_5_2 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  dirty_5_3 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  dirty_5_4 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  dirty_5_5 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  dirty_5_6 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  dirty_5_7 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  dirty_6_0 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  dirty_6_1 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  dirty_6_2 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  dirty_6_3 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  dirty_6_4 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  dirty_6_5 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  dirty_6_6 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  dirty_6_7 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  dirty_7_0 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  dirty_7_1 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  dirty_7_2 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  dirty_7_3 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  dirty_7_4 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  dirty_7_5 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  dirty_7_6 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  dirty_7_7 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  mem_rd_set_addr = _RAND_704[2:0];
  _RAND_705 = {1{`RANDOM}};
  mem_rd_tag_addr = _RAND_705[5:0];
  _RAND_706 = {1{`RANDOM}};
  mem_wr_addr = _RAND_706[8:0];
  _RAND_707 = {1{`RANDOM}};
  cacheState = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  FIFO_Choice_0 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  FIFO_Choice_1 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  FIFO_Choice_2 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  FIFO_Choice_3 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  FIFO_Choice_4 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  FIFO_Choice_5 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  FIFO_Choice_6 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  FIFO_Choice_7 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  mem_wr_line_0 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  mem_wr_line_1 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  mem_wr_line_2 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  mem_wr_line_3 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  mem_wr_line_4 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  mem_wr_line_5 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  mem_wr_line_6 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  mem_wr_line_7 = _RAND_723[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheAXI(
  input         clock,
  input         reset,
  input  [8:0]  io_mem_addr,
  input         io_mem_rd_req,
  input         io_mem_wr_req,
  input  [31:0] io_mem_wr_line_0,
  input  [31:0] io_mem_wr_line_1,
  input  [31:0] io_mem_wr_line_2,
  input  [31:0] io_mem_wr_line_3,
  input  [31:0] io_mem_wr_line_4,
  input  [31:0] io_mem_wr_line_5,
  input  [31:0] io_mem_wr_line_6,
  input  [31:0] io_mem_wr_line_7,
  output [31:0] io_mem_rd_line_0,
  output [31:0] io_mem_rd_line_1,
  output [31:0] io_mem_rd_line_2,
  output [31:0] io_mem_rd_line_3,
  output [31:0] io_mem_rd_line_4,
  output [31:0] io_mem_rd_line_5,
  output [31:0] io_mem_rd_line_6,
  output [31:0] io_mem_rd_line_7,
  output        io_cacheAXI_gnt,
  output        io_TVALID,
  output        io_TLAST,
  input         io_TREADY,
  input  [31:0] io_TDATAR,
  output [31:0] io_TDATAW,
  output [1:0]  io_TUSER
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] transferCounter; // @[CacheAXI.scala 45:32]
  reg [1:0] cacheAXIState; // @[CacheAXI.scala 47:30]
  reg  rdLine_0; // @[CacheAXI.scala 55:23]
  reg  rdLine_1; // @[CacheAXI.scala 55:23]
  reg  rdLine_2; // @[CacheAXI.scala 55:23]
  reg  rdLine_3; // @[CacheAXI.scala 55:23]
  reg  rdLine_4; // @[CacheAXI.scala 55:23]
  reg  rdLine_5; // @[CacheAXI.scala 55:23]
  reg  rdLine_6; // @[CacheAXI.scala 55:23]
  reg  rdLine_7; // @[CacheAXI.scala 55:23]
  wire [1:0] _GEN_0 = io_TREADY ? 2'h1 : cacheAXIState; // @[CacheAXI.scala 64:35 65:25 47:30]
  wire [1:0] _GEN_1 = io_mem_rd_req ? _GEN_0 : cacheAXIState; // @[CacheAXI.scala 47:30 63:37]
  wire  _T_11 = transferCounter <= 32'h8; // @[CacheAXI.scala 78:30]
  wire  _T_12 = transferCounter == 32'h0; // @[CacheAXI.scala 80:32]
  wire [31:0] _TDATAW_T = {18'h0,io_mem_addr,5'h0}; // @[Cat.scala 31:58]
  wire [31:0] _T_14 = transferCounter - 32'h1; // @[CacheAXI.scala 83:35]
  wire  _GEN_4 = 3'h0 == _T_14[2:0] ? io_TDATAR[0] : rdLine_0; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_5 = 3'h1 == _T_14[2:0] ? io_TDATAR[0] : rdLine_1; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_6 = 3'h2 == _T_14[2:0] ? io_TDATAR[0] : rdLine_2; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_7 = 3'h3 == _T_14[2:0] ? io_TDATAR[0] : rdLine_3; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_8 = 3'h4 == _T_14[2:0] ? io_TDATAR[0] : rdLine_4; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_9 = 3'h5 == _T_14[2:0] ? io_TDATAR[0] : rdLine_5; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_10 = 3'h6 == _T_14[2:0] ? io_TDATAR[0] : rdLine_6; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire  _GEN_11 = 3'h7 == _T_14[2:0] ? io_TDATAR[0] : rdLine_7; // @[CacheAXI.scala 55:23 83:{41,41}]
  wire [31:0] _GEN_12 = transferCounter == 32'h0 ? _TDATAW_T : 32'h0; // @[CacheAXI.scala 80:40 81:20]
  wire  _GEN_13 = transferCounter == 32'h0 ? rdLine_0 : _GEN_4; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_14 = transferCounter == 32'h0 ? rdLine_1 : _GEN_5; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_15 = transferCounter == 32'h0 ? rdLine_2 : _GEN_6; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_16 = transferCounter == 32'h0 ? rdLine_3 : _GEN_7; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_17 = transferCounter == 32'h0 ? rdLine_4 : _GEN_8; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_18 = transferCounter == 32'h0 ? rdLine_5 : _GEN_9; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_19 = transferCounter == 32'h0 ? rdLine_6 : _GEN_10; // @[CacheAXI.scala 55:23 80:40]
  wire  _GEN_20 = transferCounter == 32'h0 ? rdLine_7 : _GEN_11; // @[CacheAXI.scala 55:23 80:40]
  wire [31:0] _transferCounter_T_1 = transferCounter + 32'h1; // @[CacheAXI.scala 85:46]
  wire [31:0] _GEN_22 = transferCounter <= 32'h8 ? _GEN_12 : 32'h0; // @[CacheAXI.scala 78:55]
  wire  _GEN_23 = transferCounter <= 32'h8 ? _GEN_13 : rdLine_0; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_24 = transferCounter <= 32'h8 ? _GEN_14 : rdLine_1; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_25 = transferCounter <= 32'h8 ? _GEN_15 : rdLine_2; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_26 = transferCounter <= 32'h8 ? _GEN_16 : rdLine_3; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_27 = transferCounter <= 32'h8 ? _GEN_17 : rdLine_4; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_28 = transferCounter <= 32'h8 ? _GEN_18 : rdLine_5; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_29 = transferCounter <= 32'h8 ? _GEN_19 : rdLine_6; // @[CacheAXI.scala 55:23 78:55]
  wire  _GEN_30 = transferCounter <= 32'h8 ? _GEN_20 : rdLine_7; // @[CacheAXI.scala 55:23 78:55]
  wire [31:0] _GEN_31 = transferCounter <= 32'h8 ? _transferCounter_T_1 : transferCounter; // @[CacheAXI.scala 78:55 85:27 45:32]
  wire  _GEN_32 = transferCounter <= 32'h8 ? 1'h0 : 1'h1; // @[CacheAXI.scala 78:55 88:17]
  wire [1:0] _GEN_33 = transferCounter <= 32'h8 ? cacheAXIState : 2'h3; // @[CacheAXI.scala 47:30 78:55 89:25]
  wire  _GEN_34 = io_TREADY & _T_11; // @[CacheAXI.scala 77:33]
  wire [31:0] _GEN_35 = io_TREADY ? _GEN_22 : 32'h0; // @[CacheAXI.scala 77:33]
  wire [31:0] _GEN_44 = io_TREADY ? _GEN_31 : transferCounter; // @[CacheAXI.scala 45:32 77:33]
  wire  _GEN_45 = io_TREADY & _GEN_32; // @[CacheAXI.scala 77:33]
  wire [1:0] _GEN_46 = io_TREADY ? _GEN_33 : cacheAXIState; // @[CacheAXI.scala 47:30 77:33]
  wire [31:0] _GEN_48 = 3'h1 == _T_14[2:0] ? io_mem_wr_line_1 : io_mem_wr_line_0; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_49 = 3'h2 == _T_14[2:0] ? io_mem_wr_line_2 : _GEN_48; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_50 = 3'h3 == _T_14[2:0] ? io_mem_wr_line_3 : _GEN_49; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_51 = 3'h4 == _T_14[2:0] ? io_mem_wr_line_4 : _GEN_50; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_52 = 3'h5 == _T_14[2:0] ? io_mem_wr_line_5 : _GEN_51; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_53 = 3'h6 == _T_14[2:0] ? io_mem_wr_line_6 : _GEN_52; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_54 = 3'h7 == _T_14[2:0] ? io_mem_wr_line_7 : _GEN_53; // @[CacheAXI.scala 103:{20,20}]
  wire [31:0] _GEN_55 = _T_12 ? _TDATAW_T : _GEN_54; // @[CacheAXI.scala 100:40 101:20 103:20]
  wire [31:0] _GEN_57 = _T_11 ? _GEN_55 : 32'h0; // @[CacheAXI.scala 98:54]
  wire [31:0] _GEN_62 = io_TREADY ? _GEN_57 : 32'h0; // @[CacheAXI.scala 97:33]
  wire [1:0] _GEN_66 = 2'h3 == cacheAXIState ? 2'h0 : cacheAXIState; // @[CacheAXI.scala 115:21 57:24 47:30]
  wire [1:0] _GEN_67 = 2'h2 == cacheAXIState ? 2'h2 : 2'h0; // @[CacheAXI.scala 57:24 96:13]
  wire [31:0] _GEN_69 = 2'h2 == cacheAXIState ? _GEN_62 : 32'h0; // @[CacheAXI.scala 57:24]
  wire [1:0] _GEN_73 = 2'h1 == cacheAXIState ? 2'h1 : _GEN_67; // @[CacheAXI.scala 57:24 76:13]
  wire  _GEN_74 = 2'h1 == cacheAXIState ? _GEN_34 : 2'h2 == cacheAXIState & _GEN_34; // @[CacheAXI.scala 57:24]
  wire [31:0] _GEN_75 = 2'h1 == cacheAXIState ? _GEN_35 : _GEN_69; // @[CacheAXI.scala 57:24]
  wire  _GEN_85 = 2'h1 == cacheAXIState ? _GEN_45 : 2'h2 == cacheAXIState & _GEN_45; // @[CacheAXI.scala 57:24]
  assign io_mem_rd_line_0 = {{31'd0}, rdLine_0}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_1 = {{31'd0}, rdLine_1}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_2 = {{31'd0}, rdLine_2}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_3 = {{31'd0}, rdLine_3}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_4 = {{31'd0}, rdLine_4}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_5 = {{31'd0}, rdLine_5}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_6 = {{31'd0}, rdLine_6}; // @[CacheAXI.scala 123:18]
  assign io_mem_rd_line_7 = {{31'd0}, rdLine_7}; // @[CacheAXI.scala 123:18]
  assign io_cacheAXI_gnt = cacheAXIState == 2'h3; // @[CacheAXI.scala 124:40]
  assign io_TVALID = 2'h0 == cacheAXIState ? 1'h0 : _GEN_74; // @[CacheAXI.scala 57:24 59:14]
  assign io_TLAST = 2'h0 == cacheAXIState ? 1'h0 : _GEN_85; // @[CacheAXI.scala 57:24 60:13]
  assign io_TDATAW = 2'h0 == cacheAXIState ? 32'h0 : _GEN_75; // @[CacheAXI.scala 57:24]
  assign io_TUSER = 2'h0 == cacheAXIState ? 2'h0 : _GEN_73; // @[CacheAXI.scala 57:24 62:13]
  always @(posedge clock) begin
    if (reset) begin // @[CacheAXI.scala 45:32]
      transferCounter <= 32'h0; // @[CacheAXI.scala 45:32]
    end else if (2'h0 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
      transferCounter <= 32'h0; // @[CacheAXI.scala 61:23]
    end else if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
      transferCounter <= _GEN_44;
    end else if (2'h2 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
      transferCounter <= _GEN_44;
    end
    if (reset) begin // @[CacheAXI.scala 47:30]
      cacheAXIState <= 2'h0; // @[CacheAXI.scala 47:30]
    end else if (2'h0 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
      if (io_mem_wr_req) begin // @[CacheAXI.scala 68:37]
        if (io_TREADY) begin // @[CacheAXI.scala 69:35]
          cacheAXIState <= 2'h2; // @[CacheAXI.scala 70:25]
        end else begin
          cacheAXIState <= _GEN_1;
        end
      end else begin
        cacheAXIState <= _GEN_1;
      end
    end else if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
      cacheAXIState <= _GEN_46;
    end else if (2'h2 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
      cacheAXIState <= _GEN_46;
    end else begin
      cacheAXIState <= _GEN_66;
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_0 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_0 <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_1 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_1 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_2 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_2 <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_3 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_3 <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_4 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_4 <= _GEN_27;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_5 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_5 <= _GEN_28;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_6 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_6 <= _GEN_29;
        end
      end
    end
    if (reset) begin // @[CacheAXI.scala 55:23]
      rdLine_7 <= 1'h0; // @[CacheAXI.scala 55:23]
    end else if (!(2'h0 == cacheAXIState)) begin // @[CacheAXI.scala 57:24]
      if (2'h1 == cacheAXIState) begin // @[CacheAXI.scala 57:24]
        if (io_TREADY) begin // @[CacheAXI.scala 77:33]
          rdLine_7 <= _GEN_30;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  transferCounter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cacheAXIState = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rdLine_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  rdLine_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rdLine_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  rdLine_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  rdLine_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  rdLine_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  rdLine_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rdLine_7 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory(
  input         clock,
  input         reset,
  input         io_TVALID,
  input  [31:0] io_TDATAW,
  output [31:0] io_TDATAR,
  input         io_TLAST,
  input  [1:0]  io_TUSER,
  input  [11:0] io_debugMemAddr,
  output [31:0] io_debugMemData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:8191]; // @[Memory.scala 33:24]
  wire  mem_TDATAR_MPORT_en; // @[Memory.scala 33:24]
  wire [12:0] mem_TDATAR_MPORT_addr; // @[Memory.scala 33:24]
  wire [31:0] mem_TDATAR_MPORT_data; // @[Memory.scala 33:24]
  wire  mem_io_debugMemData_MPORT_en; // @[Memory.scala 33:24]
  wire [12:0] mem_io_debugMemData_MPORT_addr; // @[Memory.scala 33:24]
  wire [31:0] mem_io_debugMemData_MPORT_data; // @[Memory.scala 33:24]
  wire [31:0] mem_MPORT_data; // @[Memory.scala 33:24]
  wire [12:0] mem_MPORT_addr; // @[Memory.scala 33:24]
  wire  mem_MPORT_mask; // @[Memory.scala 33:24]
  wire  mem_MPORT_en; // @[Memory.scala 33:24]
  reg  mem_TDATAR_MPORT_en_pipe_0;
  reg [12:0] mem_TDATAR_MPORT_addr_pipe_0;
  reg  mem_io_debugMemData_MPORT_en_pipe_0;
  reg [12:0] mem_io_debugMemData_MPORT_addr_pipe_0;
  reg [1:0] memState; // @[Memory.scala 38:25]
  reg [31:0] transferCounter; // @[Memory.scala 42:32]
  reg [29:0] rwmemAddr; // @[Memory.scala 43:26]
  wire  _T_2 = 2'h0 == memState; // @[Memory.scala 45:19]
  wire [1:0] _GEN_0 = io_TUSER == 2'h2 ? 2'h2 : memState; // @[Memory.scala 51:54 52:20 38:25]
  wire  _GEN_8 = transferCounter == 32'h0 ? 1'h0 : 1'h1; // @[Memory.scala 33:24 59:38]
  wire [31:0] _GEN_11 = transferCounter == 32'h0 ? 32'h0 : mem_TDATAR_MPORT_data; // @[Memory.scala 59:38 62:18]
  wire [29:0] _rwmemAddr_T_2 = rwmemAddr + 30'h1; // @[Memory.scala 64:32]
  wire [31:0] _transferCounter_T_1 = transferCounter + 32'h1; // @[Memory.scala 65:44]
  wire [29:0] _GEN_12 = ~io_TLAST ? _rwmemAddr_T_2 : rwmemAddr; // @[Memory.scala 57:34 64:19 43:26]
  wire  _GEN_13 = ~io_TLAST & _GEN_8; // @[Memory.scala 33:24 57:34]
  wire [31:0] _GEN_16 = ~io_TLAST ? _GEN_11 : 32'h0; // @[Memory.scala 57:34]
  wire [31:0] _GEN_17 = ~io_TLAST ? _transferCounter_T_1 : transferCounter; // @[Memory.scala 57:34 65:25 42:32]
  wire [1:0] _GEN_18 = ~io_TLAST ? memState : 2'h0; // @[Memory.scala 38:25 57:34 67:18]
  wire  _GEN_42 = 2'h1 == memState & _GEN_13; // @[Memory.scala 45:19 33:24]
  wire [31:0] _GEN_45 = 2'h1 == memState ? _GEN_16 : 32'h0; // @[Memory.scala 45:19]
  wire  _GEN_50 = 2'h1 == memState ? 1'h0 : 2'h2 == memState & _GEN_13; // @[Memory.scala 45:19 33:24]
  assign mem_TDATAR_MPORT_en = mem_TDATAR_MPORT_en_pipe_0;
  assign mem_TDATAR_MPORT_addr = mem_TDATAR_MPORT_addr_pipe_0;
  assign mem_TDATAR_MPORT_data = mem[mem_TDATAR_MPORT_addr]; // @[Memory.scala 33:24]
  assign mem_io_debugMemData_MPORT_en = mem_io_debugMemData_MPORT_en_pipe_0;
  assign mem_io_debugMemData_MPORT_addr = mem_io_debugMemData_MPORT_addr_pipe_0;
  assign mem_io_debugMemData_MPORT_data = mem[mem_io_debugMemData_MPORT_addr]; // @[Memory.scala 33:24]
  assign mem_MPORT_data = io_TDATAW;
  assign mem_MPORT_addr = rwmemAddr[12:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = _T_2 ? 1'h0 : _GEN_50;
  assign io_TDATAR = 2'h0 == memState ? 32'h0 : _GEN_45; // @[Memory.scala 45:19]
  assign io_debugMemData = mem_io_debugMemData_MPORT_data; // @[Memory.scala 93:19]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 33:24]
    end
    if (_T_2) begin
      mem_TDATAR_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      mem_TDATAR_MPORT_en_pipe_0 <= _GEN_42;
    end
    if (_T_2 ? 1'h0 : _GEN_42) begin
      mem_TDATAR_MPORT_addr_pipe_0 <= rwmemAddr[12:0];
    end
    mem_io_debugMemData_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_io_debugMemData_MPORT_addr_pipe_0 <= {{1'd0}, io_debugMemAddr};
    end
    if (reset) begin // @[Memory.scala 38:25]
      memState <= 2'h0; // @[Memory.scala 38:25]
    end else if (2'h0 == memState) begin // @[Memory.scala 45:19]
      if (io_TVALID) begin // @[Memory.scala 48:33]
        if (io_TUSER == 2'h1) begin // @[Memory.scala 49:47]
          memState <= 2'h1; // @[Memory.scala 50:20]
        end else begin
          memState <= _GEN_0;
        end
      end
    end else if (2'h1 == memState) begin // @[Memory.scala 45:19]
      memState <= _GEN_18;
    end else if (2'h2 == memState) begin // @[Memory.scala 45:19]
      memState <= _GEN_18;
    end
    if (reset) begin // @[Memory.scala 42:32]
      transferCounter <= 32'h0; // @[Memory.scala 42:32]
    end else if (2'h0 == memState) begin // @[Memory.scala 45:19]
      transferCounter <= 32'h0; // @[Memory.scala 47:23]
    end else if (2'h1 == memState) begin // @[Memory.scala 45:19]
      transferCounter <= _GEN_17;
    end else if (2'h2 == memState) begin // @[Memory.scala 45:19]
      transferCounter <= _GEN_17;
    end
    if (reset) begin // @[Memory.scala 43:26]
      rwmemAddr <= 30'h0; // @[Memory.scala 43:26]
    end else if (!(2'h0 == memState)) begin // @[Memory.scala 45:19]
      if (2'h1 == memState) begin // @[Memory.scala 45:19]
        rwmemAddr <= _GEN_12;
      end else if (2'h2 == memState) begin // @[Memory.scala 45:19]
        rwmemAddr <= _GEN_12;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_TDATAR_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_TDATAR_MPORT_addr_pipe_0 = _RAND_2[12:0];
  _RAND_3 = {1{`RANDOM}};
  mem_io_debugMemData_MPORT_en_pipe_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  mem_io_debugMemData_MPORT_addr_pipe_0 = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  memState = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  transferCounter = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rwmemAddr = _RAND_7[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RPSTop(
  input         clock,
  input         reset,
  input         io_std_clk,
  input  [31:0] io_boot_addr_0,
  input  [31:0] io_boot_addr_1,
  input  [11:0] io_debugMemAddr,
  output [31:0] io_debugMemData
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  core_clock; // @[RPSTop.scala 27:20]
  wire  core_reset; // @[RPSTop.scala 27:20]
  wire  core_io_std_clk; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_boot_addr_0; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_boot_addr_1; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_instr_addr; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_instr_data; // @[RPSTop.scala 27:20]
  wire  core_io_data_we; // @[RPSTop.scala 27:20]
  wire [3:0] core_io_data_be; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_data_addr; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_data_wdata; // @[RPSTop.scala 27:20]
  wire [31:0] core_io_data_rdata; // @[RPSTop.scala 27:20]
  wire  core_io_IMiss; // @[RPSTop.scala 27:20]
  wire  core_io_DMiss; // @[RPSTop.scala 27:20]
  wire  Icache_clock; // @[RPSTop.scala 28:22]
  wire  Icache_reset; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_addr; // @[RPSTop.scala 28:22]
  wire  Icache_io_r_req; // @[RPSTop.scala 28:22]
  wire  Icache_io_w_req; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_writedata; // @[RPSTop.scala 28:22]
  wire [3:0] Icache_io_writeMask; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_outdata; // @[RPSTop.scala 28:22]
  wire  Icache_io_miss; // @[RPSTop.scala 28:22]
  wire [8:0] Icache_io_mem_addr; // @[RPSTop.scala 28:22]
  wire  Icache_io_mem_rd_req; // @[RPSTop.scala 28:22]
  wire  Icache_io_mem_wr_req; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_0; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_1; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_2; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_3; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_4; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_5; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_6; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_wr_line_7; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_0; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_1; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_2; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_3; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_4; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_5; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_6; // @[RPSTop.scala 28:22]
  wire [31:0] Icache_io_mem_rd_line_7; // @[RPSTop.scala 28:22]
  wire  Icache_io_cacheAXI_gnt; // @[RPSTop.scala 28:22]
  wire  Dcache_clock; // @[RPSTop.scala 29:22]
  wire  Dcache_reset; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_addr; // @[RPSTop.scala 29:22]
  wire  Dcache_io_r_req; // @[RPSTop.scala 29:22]
  wire  Dcache_io_w_req; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_writedata; // @[RPSTop.scala 29:22]
  wire [3:0] Dcache_io_writeMask; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_outdata; // @[RPSTop.scala 29:22]
  wire  Dcache_io_miss; // @[RPSTop.scala 29:22]
  wire [8:0] Dcache_io_mem_addr; // @[RPSTop.scala 29:22]
  wire  Dcache_io_mem_rd_req; // @[RPSTop.scala 29:22]
  wire  Dcache_io_mem_wr_req; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_0; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_1; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_2; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_3; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_4; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_5; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_6; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_wr_line_7; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_0; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_1; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_2; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_3; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_4; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_5; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_6; // @[RPSTop.scala 29:22]
  wire [31:0] Dcache_io_mem_rd_line_7; // @[RPSTop.scala 29:22]
  wire  Dcache_io_cacheAXI_gnt; // @[RPSTop.scala 29:22]
  wire  IcacheAXI_clock; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_reset; // @[RPSTop.scala 30:25]
  wire [8:0] IcacheAXI_io_mem_addr; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_io_mem_rd_req; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_io_mem_wr_req; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_0; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_1; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_2; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_3; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_4; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_5; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_6; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_wr_line_7; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_0; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_1; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_2; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_3; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_4; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_5; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_6; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_mem_rd_line_7; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_io_cacheAXI_gnt; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_io_TVALID; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_io_TLAST; // @[RPSTop.scala 30:25]
  wire  IcacheAXI_io_TREADY; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_TDATAR; // @[RPSTop.scala 30:25]
  wire [31:0] IcacheAXI_io_TDATAW; // @[RPSTop.scala 30:25]
  wire [1:0] IcacheAXI_io_TUSER; // @[RPSTop.scala 30:25]
  wire  DcacheAXI_clock; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_reset; // @[RPSTop.scala 31:25]
  wire [8:0] DcacheAXI_io_mem_addr; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_io_mem_rd_req; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_io_mem_wr_req; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_0; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_1; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_2; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_3; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_4; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_5; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_6; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_wr_line_7; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_0; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_1; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_2; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_3; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_4; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_5; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_6; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_mem_rd_line_7; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_io_cacheAXI_gnt; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_io_TVALID; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_io_TLAST; // @[RPSTop.scala 31:25]
  wire  DcacheAXI_io_TREADY; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_TDATAR; // @[RPSTop.scala 31:25]
  wire [31:0] DcacheAXI_io_TDATAW; // @[RPSTop.scala 31:25]
  wire [1:0] DcacheAXI_io_TUSER; // @[RPSTop.scala 31:25]
  wire  mem_clock; // @[RPSTop.scala 32:19]
  wire  mem_reset; // @[RPSTop.scala 32:19]
  wire  mem_io_TVALID; // @[RPSTop.scala 32:19]
  wire [31:0] mem_io_TDATAW; // @[RPSTop.scala 32:19]
  wire [31:0] mem_io_TDATAR; // @[RPSTop.scala 32:19]
  wire  mem_io_TLAST; // @[RPSTop.scala 32:19]
  wire [1:0] mem_io_TUSER; // @[RPSTop.scala 32:19]
  wire [11:0] mem_io_debugMemAddr; // @[RPSTop.scala 32:19]
  wire [31:0] mem_io_debugMemData; // @[RPSTop.scala 32:19]
  reg  cid; // @[RPSTop.scala 71:20]
  wire  _T = ~cid; // @[RPSTop.scala 82:12]
  wire [31:0] _GEN_0 = cid ? DcacheAXI_io_TDATAW : 32'h0; // @[RPSTop.scala 74:17 89:45 90:19]
  wire [1:0] _GEN_1 = cid ? DcacheAXI_io_TUSER : 2'h0; // @[RPSTop.scala 75:16 89:45 91:18]
  wire  _GEN_2 = cid & DcacheAXI_io_TVALID; // @[RPSTop.scala 76:17 89:45 92:19]
  wire  _GEN_3 = cid & DcacheAXI_io_TLAST; // @[RPSTop.scala 77:16 89:45 93:18]
  wire [31:0] _GEN_5 = cid ? mem_io_TDATAR : 32'h0; // @[RPSTop.scala 81:23 89:45 95:25]
  wire  _GEN_14 = IcacheAXI_io_TUSER != 2'h0 | cid; // @[RPSTop.scala 100:11 71:20 99:50]
  rpu_core core ( // @[RPSTop.scala 27:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_std_clk(core_io_std_clk),
    .io_boot_addr_0(core_io_boot_addr_0),
    .io_boot_addr_1(core_io_boot_addr_1),
    .io_instr_addr(core_io_instr_addr),
    .io_instr_data(core_io_instr_data),
    .io_data_we(core_io_data_we),
    .io_data_be(core_io_data_be),
    .io_data_addr(core_io_data_addr),
    .io_data_wdata(core_io_data_wdata),
    .io_data_rdata(core_io_data_rdata),
    .io_IMiss(core_io_IMiss),
    .io_DMiss(core_io_DMiss)
  );
  Cache Icache ( // @[RPSTop.scala 28:22]
    .clock(Icache_clock),
    .reset(Icache_reset),
    .io_addr(Icache_io_addr),
    .io_r_req(Icache_io_r_req),
    .io_w_req(Icache_io_w_req),
    .io_writedata(Icache_io_writedata),
    .io_writeMask(Icache_io_writeMask),
    .io_outdata(Icache_io_outdata),
    .io_miss(Icache_io_miss),
    .io_mem_addr(Icache_io_mem_addr),
    .io_mem_rd_req(Icache_io_mem_rd_req),
    .io_mem_wr_req(Icache_io_mem_wr_req),
    .io_mem_wr_line_0(Icache_io_mem_wr_line_0),
    .io_mem_wr_line_1(Icache_io_mem_wr_line_1),
    .io_mem_wr_line_2(Icache_io_mem_wr_line_2),
    .io_mem_wr_line_3(Icache_io_mem_wr_line_3),
    .io_mem_wr_line_4(Icache_io_mem_wr_line_4),
    .io_mem_wr_line_5(Icache_io_mem_wr_line_5),
    .io_mem_wr_line_6(Icache_io_mem_wr_line_6),
    .io_mem_wr_line_7(Icache_io_mem_wr_line_7),
    .io_mem_rd_line_0(Icache_io_mem_rd_line_0),
    .io_mem_rd_line_1(Icache_io_mem_rd_line_1),
    .io_mem_rd_line_2(Icache_io_mem_rd_line_2),
    .io_mem_rd_line_3(Icache_io_mem_rd_line_3),
    .io_mem_rd_line_4(Icache_io_mem_rd_line_4),
    .io_mem_rd_line_5(Icache_io_mem_rd_line_5),
    .io_mem_rd_line_6(Icache_io_mem_rd_line_6),
    .io_mem_rd_line_7(Icache_io_mem_rd_line_7),
    .io_cacheAXI_gnt(Icache_io_cacheAXI_gnt)
  );
  Cache Dcache ( // @[RPSTop.scala 29:22]
    .clock(Dcache_clock),
    .reset(Dcache_reset),
    .io_addr(Dcache_io_addr),
    .io_r_req(Dcache_io_r_req),
    .io_w_req(Dcache_io_w_req),
    .io_writedata(Dcache_io_writedata),
    .io_writeMask(Dcache_io_writeMask),
    .io_outdata(Dcache_io_outdata),
    .io_miss(Dcache_io_miss),
    .io_mem_addr(Dcache_io_mem_addr),
    .io_mem_rd_req(Dcache_io_mem_rd_req),
    .io_mem_wr_req(Dcache_io_mem_wr_req),
    .io_mem_wr_line_0(Dcache_io_mem_wr_line_0),
    .io_mem_wr_line_1(Dcache_io_mem_wr_line_1),
    .io_mem_wr_line_2(Dcache_io_mem_wr_line_2),
    .io_mem_wr_line_3(Dcache_io_mem_wr_line_3),
    .io_mem_wr_line_4(Dcache_io_mem_wr_line_4),
    .io_mem_wr_line_5(Dcache_io_mem_wr_line_5),
    .io_mem_wr_line_6(Dcache_io_mem_wr_line_6),
    .io_mem_wr_line_7(Dcache_io_mem_wr_line_7),
    .io_mem_rd_line_0(Dcache_io_mem_rd_line_0),
    .io_mem_rd_line_1(Dcache_io_mem_rd_line_1),
    .io_mem_rd_line_2(Dcache_io_mem_rd_line_2),
    .io_mem_rd_line_3(Dcache_io_mem_rd_line_3),
    .io_mem_rd_line_4(Dcache_io_mem_rd_line_4),
    .io_mem_rd_line_5(Dcache_io_mem_rd_line_5),
    .io_mem_rd_line_6(Dcache_io_mem_rd_line_6),
    .io_mem_rd_line_7(Dcache_io_mem_rd_line_7),
    .io_cacheAXI_gnt(Dcache_io_cacheAXI_gnt)
  );
  CacheAXI IcacheAXI ( // @[RPSTop.scala 30:25]
    .clock(IcacheAXI_clock),
    .reset(IcacheAXI_reset),
    .io_mem_addr(IcacheAXI_io_mem_addr),
    .io_mem_rd_req(IcacheAXI_io_mem_rd_req),
    .io_mem_wr_req(IcacheAXI_io_mem_wr_req),
    .io_mem_wr_line_0(IcacheAXI_io_mem_wr_line_0),
    .io_mem_wr_line_1(IcacheAXI_io_mem_wr_line_1),
    .io_mem_wr_line_2(IcacheAXI_io_mem_wr_line_2),
    .io_mem_wr_line_3(IcacheAXI_io_mem_wr_line_3),
    .io_mem_wr_line_4(IcacheAXI_io_mem_wr_line_4),
    .io_mem_wr_line_5(IcacheAXI_io_mem_wr_line_5),
    .io_mem_wr_line_6(IcacheAXI_io_mem_wr_line_6),
    .io_mem_wr_line_7(IcacheAXI_io_mem_wr_line_7),
    .io_mem_rd_line_0(IcacheAXI_io_mem_rd_line_0),
    .io_mem_rd_line_1(IcacheAXI_io_mem_rd_line_1),
    .io_mem_rd_line_2(IcacheAXI_io_mem_rd_line_2),
    .io_mem_rd_line_3(IcacheAXI_io_mem_rd_line_3),
    .io_mem_rd_line_4(IcacheAXI_io_mem_rd_line_4),
    .io_mem_rd_line_5(IcacheAXI_io_mem_rd_line_5),
    .io_mem_rd_line_6(IcacheAXI_io_mem_rd_line_6),
    .io_mem_rd_line_7(IcacheAXI_io_mem_rd_line_7),
    .io_cacheAXI_gnt(IcacheAXI_io_cacheAXI_gnt),
    .io_TVALID(IcacheAXI_io_TVALID),
    .io_TLAST(IcacheAXI_io_TLAST),
    .io_TREADY(IcacheAXI_io_TREADY),
    .io_TDATAR(IcacheAXI_io_TDATAR),
    .io_TDATAW(IcacheAXI_io_TDATAW),
    .io_TUSER(IcacheAXI_io_TUSER)
  );
  CacheAXI DcacheAXI ( // @[RPSTop.scala 31:25]
    .clock(DcacheAXI_clock),
    .reset(DcacheAXI_reset),
    .io_mem_addr(DcacheAXI_io_mem_addr),
    .io_mem_rd_req(DcacheAXI_io_mem_rd_req),
    .io_mem_wr_req(DcacheAXI_io_mem_wr_req),
    .io_mem_wr_line_0(DcacheAXI_io_mem_wr_line_0),
    .io_mem_wr_line_1(DcacheAXI_io_mem_wr_line_1),
    .io_mem_wr_line_2(DcacheAXI_io_mem_wr_line_2),
    .io_mem_wr_line_3(DcacheAXI_io_mem_wr_line_3),
    .io_mem_wr_line_4(DcacheAXI_io_mem_wr_line_4),
    .io_mem_wr_line_5(DcacheAXI_io_mem_wr_line_5),
    .io_mem_wr_line_6(DcacheAXI_io_mem_wr_line_6),
    .io_mem_wr_line_7(DcacheAXI_io_mem_wr_line_7),
    .io_mem_rd_line_0(DcacheAXI_io_mem_rd_line_0),
    .io_mem_rd_line_1(DcacheAXI_io_mem_rd_line_1),
    .io_mem_rd_line_2(DcacheAXI_io_mem_rd_line_2),
    .io_mem_rd_line_3(DcacheAXI_io_mem_rd_line_3),
    .io_mem_rd_line_4(DcacheAXI_io_mem_rd_line_4),
    .io_mem_rd_line_5(DcacheAXI_io_mem_rd_line_5),
    .io_mem_rd_line_6(DcacheAXI_io_mem_rd_line_6),
    .io_mem_rd_line_7(DcacheAXI_io_mem_rd_line_7),
    .io_cacheAXI_gnt(DcacheAXI_io_cacheAXI_gnt),
    .io_TVALID(DcacheAXI_io_TVALID),
    .io_TLAST(DcacheAXI_io_TLAST),
    .io_TREADY(DcacheAXI_io_TREADY),
    .io_TDATAR(DcacheAXI_io_TDATAR),
    .io_TDATAW(DcacheAXI_io_TDATAW),
    .io_TUSER(DcacheAXI_io_TUSER)
  );
  Memory mem ( // @[RPSTop.scala 32:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_TVALID(mem_io_TVALID),
    .io_TDATAW(mem_io_TDATAW),
    .io_TDATAR(mem_io_TDATAR),
    .io_TLAST(mem_io_TLAST),
    .io_TUSER(mem_io_TUSER),
    .io_debugMemAddr(mem_io_debugMemAddr),
    .io_debugMemData(mem_io_debugMemData)
  );
  assign io_debugMemData = mem_io_debugMemData; // @[RPSTop.scala 110:19]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_std_clk = io_std_clk; // @[RPSTop.scala 35:19]
  assign core_io_boot_addr_0 = io_boot_addr_0; // @[RPSTop.scala 36:21]
  assign core_io_boot_addr_1 = io_boot_addr_1; // @[RPSTop.scala 36:21]
  assign core_io_instr_data = Icache_io_outdata; // @[RPSTop.scala 37:22]
  assign core_io_data_rdata = Dcache_io_outdata; // @[RPSTop.scala 38:22]
  assign core_io_IMiss = Icache_io_miss; // @[RPSTop.scala 39:17]
  assign core_io_DMiss = Dcache_io_miss; // @[RPSTop.scala 40:17]
  assign Icache_clock = clock;
  assign Icache_reset = reset;
  assign Icache_io_addr = core_io_instr_addr; // @[RPSTop.scala 43:18]
  assign Icache_io_r_req = 1'h1; // @[RPSTop.scala 52:19]
  assign Icache_io_w_req = 1'h0; // @[RPSTop.scala 45:19]
  assign Icache_io_writedata = 32'h0; // @[RPSTop.scala 46:23]
  assign Icache_io_writeMask = 4'h0; // @[RPSTop.scala 44:23]
  assign Icache_io_mem_rd_line_0 = IcacheAXI_io_mem_rd_line_0; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_1 = IcacheAXI_io_mem_rd_line_1; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_2 = IcacheAXI_io_mem_rd_line_2; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_3 = IcacheAXI_io_mem_rd_line_3; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_4 = IcacheAXI_io_mem_rd_line_4; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_5 = IcacheAXI_io_mem_rd_line_5; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_6 = IcacheAXI_io_mem_rd_line_6; // @[RPSTop.scala 56:25]
  assign Icache_io_mem_rd_line_7 = IcacheAXI_io_mem_rd_line_7; // @[RPSTop.scala 56:25]
  assign Icache_io_cacheAXI_gnt = IcacheAXI_io_cacheAXI_gnt; // @[RPSTop.scala 57:26]
  assign Dcache_clock = clock;
  assign Dcache_reset = reset;
  assign Dcache_io_addr = core_io_data_addr; // @[RPSTop.scala 47:18]
  assign Dcache_io_r_req = 1'h0; // @[RPSTop.scala 53:19]
  assign Dcache_io_w_req = core_io_data_we; // @[RPSTop.scala 49:19]
  assign Dcache_io_writedata = core_io_data_wdata; // @[RPSTop.scala 50:23]
  assign Dcache_io_writeMask = core_io_data_be; // @[RPSTop.scala 48:23]
  assign Dcache_io_mem_rd_line_0 = DcacheAXI_io_mem_rd_line_0; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_1 = DcacheAXI_io_mem_rd_line_1; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_2 = DcacheAXI_io_mem_rd_line_2; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_3 = DcacheAXI_io_mem_rd_line_3; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_4 = DcacheAXI_io_mem_rd_line_4; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_5 = DcacheAXI_io_mem_rd_line_5; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_6 = DcacheAXI_io_mem_rd_line_6; // @[RPSTop.scala 58:25]
  assign Dcache_io_mem_rd_line_7 = DcacheAXI_io_mem_rd_line_7; // @[RPSTop.scala 58:25]
  assign Dcache_io_cacheAXI_gnt = DcacheAXI_io_cacheAXI_gnt; // @[RPSTop.scala 59:26]
  assign IcacheAXI_clock = clock;
  assign IcacheAXI_reset = reset;
  assign IcacheAXI_io_mem_addr = Icache_io_mem_addr; // @[RPSTop.scala 62:25]
  assign IcacheAXI_io_mem_rd_req = Icache_io_mem_rd_req; // @[RPSTop.scala 63:27]
  assign IcacheAXI_io_mem_wr_req = Icache_io_mem_wr_req; // @[RPSTop.scala 64:27]
  assign IcacheAXI_io_mem_wr_line_0 = Icache_io_mem_wr_line_0; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_1 = Icache_io_mem_wr_line_1; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_2 = Icache_io_mem_wr_line_2; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_3 = Icache_io_mem_wr_line_3; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_4 = Icache_io_mem_wr_line_4; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_5 = Icache_io_mem_wr_line_5; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_6 = Icache_io_mem_wr_line_6; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_mem_wr_line_7 = Icache_io_mem_wr_line_7; // @[RPSTop.scala 65:28]
  assign IcacheAXI_io_TREADY = ~cid; // @[RPSTop.scala 82:12]
  assign IcacheAXI_io_TDATAR = ~cid ? mem_io_TDATAR : 32'h0; // @[RPSTop.scala 79:23 82:39 88:25]
  assign DcacheAXI_clock = clock;
  assign DcacheAXI_reset = reset;
  assign DcacheAXI_io_mem_addr = Dcache_io_mem_addr; // @[RPSTop.scala 66:25]
  assign DcacheAXI_io_mem_rd_req = Dcache_io_mem_rd_req; // @[RPSTop.scala 67:27]
  assign DcacheAXI_io_mem_wr_req = Dcache_io_mem_wr_req; // @[RPSTop.scala 68:27]
  assign DcacheAXI_io_mem_wr_line_0 = Dcache_io_mem_wr_line_0; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_1 = Dcache_io_mem_wr_line_1; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_2 = Dcache_io_mem_wr_line_2; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_3 = Dcache_io_mem_wr_line_3; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_4 = Dcache_io_mem_wr_line_4; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_5 = Dcache_io_mem_wr_line_5; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_6 = Dcache_io_mem_wr_line_6; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_mem_wr_line_7 = Dcache_io_mem_wr_line_7; // @[RPSTop.scala 69:28]
  assign DcacheAXI_io_TREADY = ~cid ? 1'h0 : cid; // @[RPSTop.scala 80:23 82:39]
  assign DcacheAXI_io_TDATAR = ~cid ? 32'h0 : _GEN_5; // @[RPSTop.scala 81:23 82:39]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_TVALID = ~cid ? IcacheAXI_io_TVALID : _GEN_2; // @[RPSTop.scala 82:39 85:19]
  assign mem_io_TDATAW = ~cid ? IcacheAXI_io_TDATAW : _GEN_0; // @[RPSTop.scala 82:39 83:19]
  assign mem_io_TLAST = ~cid ? IcacheAXI_io_TLAST : _GEN_3; // @[RPSTop.scala 82:39 86:18]
  assign mem_io_TUSER = ~cid ? IcacheAXI_io_TUSER : _GEN_1; // @[RPSTop.scala 82:39 84:18]
  assign mem_io_debugMemAddr = io_debugMemAddr; // @[RPSTop.scala 109:23]
  always @(posedge clock) begin
    if (reset) begin // @[RPSTop.scala 71:20]
      cid <= 1'h0; // @[RPSTop.scala 71:20]
    end else if (_T) begin // @[RPSTop.scala 98:39]
      cid <= _GEN_14;
    end else if (cid) begin // @[RPSTop.scala 102:45]
      if (DcacheAXI_io_TUSER != 2'h0) begin // @[RPSTop.scala 103:50]
        cid <= 1'h0; // @[RPSTop.scala 104:11]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cid = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
